�P  ��> @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �              �      p     �             �            �             �             <      �      ?�      �      {�@     �      �@     �     w�      �     �      �      ���     �      ���     �      o��     �      ��    ��      /��     �      ?��    ��      ��     �      ��    ��      ��     �      ��    ��      8?      �      ?�     ��      <      �      ?�     À      >>      �      ?�     ��      |              |      �      (:              (:      �      @               @       �                              �                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        > > �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ������� ������� ������� ������� ������� ������� ������� ������  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  ������  ������  ������  ������  ������  ������  ������  ������@������@������@������@�������������������������������������������������������������������������������������������?�������?�������?�������?���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �   � � �   � � �   � � �   � � �                                > @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            8       8       8                               �       �             �     �      �       >      �     �>      �       >�     ��    �>�     ��      >      ��    �>     �          ��    �     ��     �     ��     ��     ���     ��    ���     �     ���     ��    ���    p�     ���     ��    ���    ��     ���     ��    ���    ��   ���    ��   ���   ��     ���     ��    ���    p��    ���     ���    ���    ���    ���    ���    ���    	���    ���    ���    ���    ���    ���    ��     ���    ��     ���    ��     ���    ��     ��     ��     ��     ��      ��     ��     ��     ��            �     �       �     ��      ��     ��       x      ��      ��      ��             ��      ��      ��               @             @             ~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            > > ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ������ ������ ������ ������  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  ?�����  ?�����  ?�����  ?�����  �����  �����  �����  �����  �����  �����  �����  ����   ����   ����   ����   ����   
����   
����   
����   
����   ����   ����   ����   �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  ?�����  ?�����  ?�����  ?�����  �����  �����  �����  �����  �����  �����  �����  �����  ������  ������  ������  ������ ������ ������ ������ ���������������������������������� ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  � � �   � � �                                                     ` > @                                                                                                                                                                                                                                                                                                                                                                              �             �             � @           � @           <�    �     ?��    �     x      �    �     �    ��       �    ���     ��     �     @�     @��    @��    ��     ?�     !��     ?��    ��     ?�     ��    8?��    ��?�    ?�     ��?�   |?��    ���    ?�     ���   |?��    ����    ?�     ����   ~?�      ��     �     ���   ���     ���     �      ���   ��     {��     u�    }ǜ   ���    ���     ��    ���   ���    ����    ���    ����  ���    ����    ����   ����   q����   ����    ���   ���   �����   �����   ����   �����   ���� 
������ 
��� 
������� 
?��  �����   ��   ����   ���   �����   ?��   ?����   ���   ����    ?��    ?���   ���    ����    ?��    ?���   ���    ����    ?��    ?���   ���    ���<@   ?���   ?���@   ����   ���    ���   ���    ����   ���    �;�   ��?�    ?���   ���    �3�   ��?�    ���   ��0�   �9�   ��?��   ���    ���     �      ��c�     ��      �     ��     ��     ��     |     }     }|    r�     |            |     ��    @|           @|    ��    �8            �8    ��                        �                              �          @               @   �                               �                                                                                                                                                                                                                                                                                                                                                                                                            > > ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?�������?�������?�������?����������������������������������������������������������� ~������ ~������ ~������ ~����}  =����}  =����}  =����}  =�����  �����  �����  �����  �����   �����   �����   �����   �����   �����   �����   �����   �����   ����   ����   ����   ����   ����   ����   ����   ����   o����   o����   o����   o���   ����   ����   ����   ����   ����   ����   ����   ����  c����  c����  c����  c����   ����   ����   ����   ����<   ���<   ���<   ���<   ����   ?����   ?����   ?����   ?���    ���    ���    ���    ���    ���    ���    ���    ��@     \�@     \�@     \�@     \��    ?���    ?���    ?���    ?���    ���    ���    ���    ���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����  ���  ���  ���  ��� ���� ���� ���� ����� F?����� F?����� F?����� F?��������������������� ������ ������ ������ �����������������������������|�=����|�=����|�=����|�=��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                        > @                                                                     �               �                                               �               �                  �               �                    �       �       �             �       �     �       >    �     �>     �                �           B         B            ���    ���    ���           ����   ����   ����     <    ����   ﻟ�  
 ����        >?��  >?�� >?��         �_�   ��   �_�    p     ���~�   ��~_� ���~_�    � @   �����  �� ��  ������   � �   q����  ����� ������   ���   �����  9����� ������  8���  �w���  }����� ������  |����  ������  }����� ������  | ��  �����߀ |����������߀ | ��   ��?��?� 8������ ������� 8 ���� p���?� ����?�w����?� ���    ����� ����� ����� ����   !������ ������ ?������ ����  A�����p ?������ ������ ?����?�A�����p ?������������ ?�����  �����0X+������x������X+������ ����0 ������?������ ������ �����0 ������������ �����������` ����������� �����������@ ������������� ����?� ����� ����� ����� ����  ������  �����  ������  ����  �����0  ?����� ������  �����  �����  ?�����  ������  �����  ?���ߜ  ?���/�  ?�����  ���#�  ?����  ?���s�  ?�����  ���s�  ?����<  ?��1�  ?�����  ��!�  �����  ?��   ?�����   ��    �����@ �?���  �����@  |?��   ������ ����  ������   ��   ����@ ����  �����@  ��    �'��  G��  �?��   @�@   ����  ���  ����   �   !�����  @����  a�����  @��  C�����   ����  C�����   ��   �����   �����  ������   ���  w?���   �?�� �?���   � �  ����   ���� ����   � �   �����  ����  �����  � �   ����@  ����  ����@  � �   ����   p~���  ����   p �   ���     ��   ���      �   �?�      ?~    �?�            �?�      ?�    �?�              �      �      �              �      �      �              �      �      �                                                                                                                   > > ���������������������������������������������������������������������������������������������������������������������������������������������������������������|�������|�������|�������|����������������������������������������������������������������������������������������������������������������������������������������������� `����� `����� `����� `����� @@���� @@���� @@���� @@���� @`���� @`���� @`���� @`������@������@������@������@���� ����� ����� ����� ��� ���� ���� ���� ����.   ��.   ��.   ��.   ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     |�     |�     |�     |�    @<�    @<�    @<�    @<�    ��    ��    ��    ���  ���  ���  ���  ���   ��   ��   ��   ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     ��     ��     ��     ��    ��    ��    ��    ��     ��     ��     ��     �x     <�x     <�x     <�x     <��    |��    |��    |��    |�`    ��`    ��`    ��`    ��     ��     ��     ��     ��@    ��@    ��@    ��@    ���    ���    ���    ���    ���   ���   ���   ���   ���   
���   
���   
���   
���    ���    ���    ���    ���    ���    ���    ���    ���    ��    ��    ��    ��  ` ���  ` ���  ` ���  ` ���� � ���� � ���� � ���� � ����   ����   ����   ����   ���    ���    ���    ���    ���    ���    ���    ���    ��x @   ��x @   ��x @   ��x @   ��� �  ��� �  ��� �  ��� �  ����  ����  ����  ����  ����  |���  |���  |���  |���  ����  ����  ����  ����  ?����  ?����  ?����  ?����  �����  �����  �����  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                        > @                                                                     �      �       �                                              �       �       �                @�       �     @�            �       �       �              �     �    �           �>   �>   �>          �    �    �            B   B   B             ���    ���    ���           ����   ����   ����          
 ����  
 ����  
 ����         >?�� >?�� >?��           �_�   �_�   �_�         ���~_� ���~_� ���~_�    |    ����  ���� ����    �    �� �� �� �� �� ��   �    �� �� �� �� �� ��   ��   �� �� �� �� �� ��   ��   �� q�� �� �� �� ��   ���  �� g�߀�� �߀�� �߀  ���   �| G�� �| ?�� �| ��  ����  v? ��?�v8 ��?�v? ��?� ��?�   ���� `��� ����  �>?�   ?������ ?�s���� ?������   |�   ������ ������ ������   ��  ������������������  ��  @������@������@������8 ��  ?�����?�����?�����| ��   ��� �� ��� �� ��� ��|  ��  �q� ����� ����� ��| ��  ��� ����� ����� �8>|���  ��  o� ��� o� ��� o� > ?���  ���> p  ���� p  ���� p  > ?��� ��� p ���� p ���� p   ���  ���x  ��� x  ����x    ���  ?���  ?�� �  ?����   ��   ?�?��  ?���  ?����   ?��>   ?���@ ?���  ?����@  ?��<   ?�_��  ?� ��  ?�_���   ��8   �����@ �  ?�@ �����@        �_���� �  ?�� �_����  �     �o���@ �` ?�@ �o���@  ?�     ���   p �  ���   ?�     ����  � ?�  ����         a�����  a�� �  a�����         C�����  C�� � C�����          ������  ������  ������   p     ?��� ?��� ?���   �     ��� ��� ���  �      ���� ���� ���� �      ���@ ���@ ���@ �      ��  ��  ��   �      ��   ��   ��    p      �?�    �?�    �?�            �?�    �?�    �?�              �     �      �             �       �       �             �      �      �                                                                                                                  > > ���������������������������������������������������������������������������������������������������������������������������������������������������������������|�������|�������|�������|��������������������������������}�������}�������}�������}������������������������������������������������������������������������������������������ `����� `����� `����� `����� @@���� @@���� @@���� @@���� @`���� @`���� @`���� @`������@������@������@������@���� ����� ����� ����� ��� ���� ���� ���� ����.  ���.  ���.  ���.  ���   ���   ���   ���   ���   `��   `��   `��   `��    ��    ��    ��    ��    ��    ��    ��    ��    |�    |�    |�    |�   @<�   @<�   @<�   @<�   ��   ��   ��   ���   ���   ���   ���   ���    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     ��     ��     ��     ��    ��    ��    ��    ��    ��    ��    ��    �@     <�@     <�@     <�@     <��    |��    |��    |��    |�@    ��@    ��@    ��@    ��     ��     ��     ��     ��@    ��@    ��@    ��@    ���    ���    ���    ���    ���    ���    ���    ���    ���   ���   ���   ���   ���    ���    ���    ���    ���    ���    ���    ���    ���    ��    ��    ��    ��    ���    ���    ���    ����   ����   ����   ����   ����   ����   ����   ����   ���    ���    ���    ���    ���    ���    ���    ���    ��x @   ��x @   ��x @   ��x @   ��� �  ��� �  ��� �  ��� �  ����  ����  ����  ����  ����  |���  |���  |���  |���  ����  ����  ����  ���� �?���� �?���� �?���� �?���� ������ ������ ������ �����������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                        > @                                                                                                                                                                                                                                                                                                                                 |       |       |              �     �     �             �     �     �      �     �      �      �       �     �      �      �       �     �      �      �       ?�    ��   ��   ��     ?�     ��    ��    ��     ?�     ��    ��    ��     ?�     ��    ��    ��     ?�     ��    ��    ��     �    ��   ��   ��     �     88   �88   �88     ��    �    ��    ��      �    >�     ?��     ?��       �    �   �  ��   �  ��   �    ��   !�     !��     !��        ��   ��     ��     ��       ��   �F     ��     ��       9��   ��     ��     ��       ���  �   8  �   8  �   8   ����  �   |  �   |  �   |   ����     ~  �  ~  �  ~   ����   �  ~   ���~   ���~   �   �  �   ����   ����  ? 8�    �  �   �� �   �� �  � �     � �   ���   ���  �� �     | �   ���   ���  �� �     ~ �   O���   O��� �� �      �   ����   ���� � �     ��?   G��?   G��? ��@�    ��    ��    ��  ���      ���    ���    ���  ��@      ���    ���    ���   ��       ���    ���    ���   ��       ���    ���    ���   � p     ���   ���   ���  ?� �     x��   x��   x��  � �    ���  ���  ���    �     ����   ����   ����     p     ?���   ?���   ?���          ���  ���  ���           ����   ����   ����           �      �      �                                                                                                                                             @       @       @                                                                                                                                                                                   > > ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ������� ������� ������� ������� ?������ ?������ ?������ ?������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������  ?�����  ?�����  ?�����  ?�����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  ����   �|��   �|��   �|��   �|��   ����   ����   ����   ����    ����    ����    ����    ����    ����    ����    ����    ����    ���    ���    ���    ���    G���    G���    G���    G���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ��     ��     ��     ��     ��     ��     ��     ��     ��     ?��     ?��     ?��     ?��     ��     ��     ��     ��     ���     ���     ���     ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ?���    ?���    ?���    ?����   ?����   ?����   ?����   ?����   |���   |���   |���   |���   �?���   �?���   �?���   �?���   ����   ����   ����   ����  ����  ����  ����  ����� ����� ����� ����� ����� �?���� �?���� �?���� �?���� ?|���� ?|���� ?|���� ?|���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                        > @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     p       p       p              |       |       |      �       �       �       �             �      �      �              �      �      �              �      �      �              �      �      �              �      �      �      >       �       �       �      >                              ��        p       p       p    ��        �       �       �    ��      �      �      �    ��>      �      �      �    ��>      �      �      �    ��>      �      �      �    ��    0 <p    0 <p    0 <p    ��     ` x     ` x     ` x     ��     � �     � �     � �           �       �       �       >      �       �       �              |�     |�     |�             8�     8�     8�              `      `      `       �      �      �      �              �      �      �              �      �      �              �      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   > > �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ������  ������  ������  ������  ������  ������  ������  ������  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  �����  ����� ����� ����� ����� ����� ������ ������ ������ ������ ������ ������ ������ ����� ������ ������ ������ ������ ������� ������� ������� �����������������������������������������������������������������?�������?�������?�������?�������������������������������������������������������������������������������������������?�������?�������?�������?�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                        > @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �      �                      �      �                      ?�      ?�                      �      �                      ��      ��                     ��      ��              �      ��      ��              �      ��      ��              �      ��      ��              �      �      �              �      ?�      ?�                     �      �                     �      �              >      ��     ��              >      ��     ��              >      ��     ��                    �8     �8                     �      �                      �      �                      ��     ��                      �      �                      �      �                      �      �                      �      �                      @       @                       �       �                       @       @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    > > ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?�������?�������?�������?�������������������������������������������������������������� ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ������ ��������������������������������������������������������������� ������� ������� ������� ������� ������� ������� ������� ������@ ������@ ������@ ������@ ��������������������������������������������������������������������������������������������������������������?�������?�������?�������?�������|������|������|������|�������?�������?�������?�������?�������?�������?�������?�������?�������?�������?�������?�������?�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                        