�P  XM' +                                                                                                                                               |    |         |    �    �         �    �    �         �   �   �        �   ��  ��        �  ��  ��        L  ?��  ?��           ��  ��       @�  ���  ���       �� � � ���    � ��� ���  �     ��� ���   |       ��� ��  @   l  �� ���  D�   8  � �}�  }�      �8 ���  }�   � �  ��� ��  D �  ���  ��  80 ? K ?��  �� >  0 ?|� ?��  � ?    �� ��  �  ?  �� ��  �  ~   ~� ~��  �� ~   |� |��  �� |   x� x��  �� x  p � p�� p�     �?�� �?�� �     0  ��� ��� �     `  ��� ��� �    
   x ~ � n �       ~ ~ �� n ��   �  < ~ � ~ � | �   � ~ � ~ p > �   $ �  � � � �  �    � �  � �  � �  8       � � � �            <      �      ?�      �   ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� O��� O��� O��� O��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��  ��  ��  ��  ��8  ��8  ��8  ��8  ��x  ��x  ��x  ��x  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ��  ��  ��  ��  � �> � �> � �> � �> ��������� ���� ���� ���� ���� ��� ��� ��� �����������������������������������������������������������������������                                    ' +                                                               >    >         >    �   �        �   ��   ��        �   ��  ��        `  ��  ��        �  �   ��   �   `  ��  ��   �   �   �  �   A    ��  �X  ��   P  ��  �  ��   �     ?�  ?��   �  0 r @� @�� @ �  `  @��?  ��� @    @�� ����  ��� �    @� ��� C��� � �  �   ��� ���� ��� �    ��� ���� ��� �    C�� ���� ��� �    �  ���� ��� �    ��  o��� ��� `   /�| ��� P�� |   ��� ���� ���  0 �� ��� ���   0 �� ��� ���   0 �� ��� ���   7 � ��� ���    ? < � <��  ��    ?  |  ��  ��    ?     ��  ��   ?   �  ��  �    ?  ?��  ?��       0   ��  ��       `   ��  ��            n   ~           ~ n  ~ ~           | ~  | ~    |       < ~  < ~    >       | �  | �  ` �        �  | �  x �  �       � ~ � ~      ������������������������������������' + �������������������������������������������������������������������������������������������������� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��   ��   ��   ��   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��8  ��8  ��8  ��8  � x  � x  � x  � x  � �  � �  � �  � �  � �  � �  � �  � �  � �  � �  � �  � �  ��  ��  ��  ��  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���> ���> ���> ���> �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������' +                                   >   ~    �   �           �  �           �   �      �� �� @    ��� ��        �  �      ? ?� ? ?�        ~� ~�    @@���� ����    
 �� ���� ����     �   ���� ����      ���������   �   ?����?����   �     ��� ���� 8 �     �� ��� ��      �� ��  �       ��  ���  ��  �    ��  ��  ��       �  ��  ��          ��  ��          ��  ��       |  ��  ��      �  ��  ��   0  ��  ��  ��    0  ��  ��  ��       ��  ��  ��    '  �  ��  ��    /   �  ��  ��    ?  |  ��  ��    ?     ��  ��   ?   �  ��  �    ?  ?��  ?��           ��  ��       @   ��  ��            ~   n           ~ ~  ~ n           | ~  | ~    |       < ~  < ~    >       | �  | �  ` �        �  | �  x �  �       � ~ � ~                                          ' + ����������������������������������������� ���� ���� ���� ����
����
����
����
��������������������?�?��?�?��?�?��?�?�����������������������������������������������������   �   �   �   �    �    �    �    �    ~    ~    ~    ~�   ~�   ~�   ~�   ~�   >�   >�   >�   >�   >�   >�   >�   >�   ~�   ~�   ~�   ~��  ���  ���  ���  ��p  ��p  ��p  ��p  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���> ���> ���> ���> �����������������������������������������������������������������������������������������������������������������������������������������  ��      ��     ��     ��     �' +                                                                                                                           |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��       ��  �  ��   �   @   �  ��  �  �0  <Dx  ?��  ��      ||  ��  ��  @l  �D�  ��  �   �8 ��� ���   |     �9� ��   �   8 �9� ���   �   8 ��� �}�   |       �ǟ ���  ��   8  ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��      �  ���  ��      �| ���  ��    �� ���  ��   ��� ���  ��   0 �� ���  �� � ? ��_ ���  �� � ? ��_ ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ������������������������������������' + �������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ���������������������������������������������������������������������������������� 
����   
����   ����   ����   ��' +                                                                                                                                               |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��       ��  �  ��   �   @   �  ��  �  �0  <Dx  ?��  ��      ||  ��  ��  @l  �D�  ��  �   �8 ��� ���   |     �9� ��   �   8 �9� ���   �   8 ��� �}�   |       �ǟ ���  ��   8  ��� ���  ��      ��� ���  ��      �� ���  ��    �  ���  ��    � / ���  ��    �|k ���  C��    =�y ���  ��     �� ���  �� �  ��_ ���  �� � ? ��_ ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ������������������������������������' + ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������  ����   ~?�      ��     �     �' +                                                                                                                                               |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��        x  ��  ��       d F  ���  ���       ��  ���  ���       �� � � ���    � ��� ���  �   A �ǿ ���   |   @ ��? ���  @  l� �� ���  D�  9  �( ���  }�   �  �8 ���  }�   � �  ���  ��  D �  ���  ��  8 �  ���  ��    � O ���  ��   0 �|� ���  �    0 ��� ���  �  �7 ��� ���  �  � ? ��_ ���  �� � ? ��_ ���  �� � ? ��_ ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �        @   �                            ' + ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ���������������������������������������������������������������������������������������������������� ~������ ~��' +                                                                                                                                                                  �   �        �   �   �            ?�   ?�        0   ��   ��        �   ?�   ��   �    0   �   ��   �    @   �� ��� �     `�  ?��  ���  �@     ?�� �� @   �� ?�� ��� �        �� ��� �        �� ��� �      �ǿ  ��  ��      �� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��   ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      �� ���� ����� F?����� F?����� ' + ������������������������������������������������������������������������������������������������������������������������������������������������������������������?����?����?����?����������������������������������� ��� ��� ��� ��� ��� ��� ��� ���  ���  ���  ���  ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������    �       �       �             ' +                                                                                                                           �    �         �   �   �        �   �   �            �   �        �   �   �        �       �   `   �   +?   ?�   �       !�   !�         5�  ?��  �   
�  @�  ��  ?�   @ F  ���  ���  #    �   ���  ���      �  �� ���      � ��� ���        �� ���   �      ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��   ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ��� ����� ����  ������  ����� ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� G��� G��� G��� G��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������                                    ' +                                                                                                                           |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��       ��  �  ��   �       �  ��  �   �   D@  ��  ��   @  p  ��  ��  l0  >D�  ?��  �    8  ��  }�|   |   @   �}�  ���   �   �  ��� �}�   |     ��� ���       8 ��� ���         ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��      �  ���  ��    �| ���  ��    �� ���  ��  0 ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ��   ��   ��   ��    ��  ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������  ?����  ?����  ?����  �����  ��' +                                                                                                                           >    >         >    �   �        �   ��   ��        �   ��  ��        `  ��  ��        �  �   ��   �   `  ��  ��   �   �   �  �   A    ��  ;�X  ;��   P  :��  ��  ���   �  �   ��  ���   �  � r �� ���   �    ��? ���       � ��� ���        �� ���   �      ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��  0 ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      �� �� �� �� ��   �    �� �� ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ���������������������������������������������������������������������������������� � ?�  ����         a�����  a��' +                                                                                                                                                                   �   �        �   �   �            �   �           ?�   ?�            �   �       @  ��  ��    
  �  ��  ��         ��  ��     `� ���� ����   � � ��������   �    ��� ����   �    ��� ��� ��    ��� ���  �       ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��  0 ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ������������������������������� ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������������?����?����?����?������������������������������������������������������������������� ��� ��� ��� ���  ���  ���  ���  ���  ~��  ~��  ~��  ~�   ~�   ~�   ~�   ~�   >�   >�   >�   >�   >�   >�   >�   >�   ~�   ~�   ~�   ~�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������  ���    ���    ���    ���    �