�3  �x ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��            ��_�                                                        �����            ��_�                                                        �����            ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �       ��_�                                                        �����     �       ��_�                                                        �����     �       ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �       ��_�                                                        �����     �       ��_�                                                        �����     �       ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �       ��_�                                                        �����     �       ��_�                                                        �����     �       ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �y͠    ��_�                                                        �����     �y͠    ��_�                                                        �����     �y͠    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �}�    ��_�                                                        �����     �}�    ��_�                                                        �����     �}�    ��_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �}�   ���_�                                                        ������   �}�   ���_�                                                        ������   �}�   ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �}�   ���_�                                                        ������   �}�   ���_�                                                        ������   �}�   ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �T"    ���_�                                                        ������   �T"    ���_�                                                        ������   �T"    ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �T�    ���_�                                                        ������   �T�    ���_�                                                        ������   �T�    ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �U"    ���_�                                                        ������   �U"    ���_�                                                        ������   �U"    ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ��     �U�    ��_�                                                        �����     �U�    ��_�                                                        �����     �U�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �U�    ��_�                                                        �����     �U�    ��_�                                                        �����     �U�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �U�    ��_�                                                        �����     �U�    ��_�                                                        �����     �U�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �T�    ��_�                                                        �����     �T�    ��_�                                                        �����     �T�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �                                                     π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �                                                     π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �                                                      �! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �                                                      �! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  ���������������������������������������������������������! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  ���������������������������������������������������������! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  ���������������������������������������������������������! ��              ��_��������������������������������������������������������������              ��_��������������������������������������������������������������              ��_������������������������������������������������������������ ��_������������  ���������������������������������������������������������! ��              ��_��������������������������������������������������������������              ��_��������������������������������������������������������������              ��_������������������������������������������������������������ ��_������������                                                            ! ��              ��_��������������������������������������������������������������              ��_��������������������������������������������������������������              ��_������������������������������������������������������������ ��_������������                                                            ! ��              ��_��������������������������������������������������������������              ��_��������������������������������������������������������������              ��_������������������������������������������������������������ ��_������������                                                            ! ��              ��_��������������������������������������������������������������              ��_��������������������������������������������������������������              ��_������������������������������������������������������������ ��_������������                                                            ! ��              ��_��������������������������������������������������������������              ��_��������������������������������������������������������������              ��_������������������������������������������������������������ �@         
�<                                                            ! ���           ���_���������������������������������������������������������������           ���_���������������������������������������������������������������           ���_������������������������������������������������������������ ������������<                                                            ! ���           ���_���������������������������������������������������������������           ���_���������������������������������������������������������������           ���_������������������������������������������������������������ �          �<                                                            ! ���           ���_���������������������������������������������������������������           ���_���������������������������������������������������������������           ���_������������������������������������������������������������ �������������<                                                            ! ���           ���_���������������������������������������������������������������           ���_���������������������������������������������������������������           ���_������������������������������������������������������������ �           �<                                                            ! ���           ���@                                                          	����           ���@                                                          	����           ���@                                                          	� �������������<  ����������������������������������������������������������� �������������������@                                                          	��������������������@                                                          	��������������������@                                                          	�                                                                               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                   @                                                          	 �������������������                                                           ��������������������                                                           ��������������������                                                           �                                                                               �������������������                                                           ��������������������                                                           ��������������������                                                           �                                                                               ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                  ������������������������������������������������������������ ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ��               �����������������������������������������������������������������               �����������������������������������������������������������������               ���������������������������������������������������������������                      8    � p        �  P      �  �  $  � �  �  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ ���������������         (  
   � @         @  P      @  �  $  �    �  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                    (  
   � @         @  P      @  �  $  �    �  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                    (      p        �  p      �  �  $  � �  �  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                    (  
             @         @  �  $  
     �  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                    (  
             @         @  �  $  
     �  ������������{��{����������������������������������������������������������������������������{��{����������������������������������������������������������������������������{��{����������������������������������������������������������������  ! ` � �         8      p        �        �  �  $  � �  �  ������������s��;����������������������������������������������������������������������������s��;����������������������������������������������������������������������������s��;����������������������������������������������������������������  c p � �                                                               ��������c��c��������������������������������������������������������������������������c��c��������������������������������������������������������������������������c��c������������������������������������������������������������������  � x� � �                                                               ��������!��C�����    �  �  p    ���  �  8    �  �  8    �  �  8    ���������!��C�����    �  �  p    ���  �  8    �  �  8    �  �  8    ���������!��C�����    �  �  p    ���  �  8    �  �  8    �  �  8    � � |� � � �����      @         �          �          �        ��� ����� �������    �  �  w������������  ;���  ����  ;���  ����  ;���  ���� ����� �������    �  �  w���������  �������  �  ����  �������  8  ������� ����� �������    �  �  w���������  �  8  ����������    �  ����������� � ~� � �        ���  ���     �          �  #������?������������ ��������!��C�����    �  �  w������������  ;���  ����  ;���  ����  ;���  ���������!��C�����    �  �  w���������  �������  �  ����  �������  8  ������������!��C�����    �  �  w���������  �  8  ����������    �  ����������� � |� � �        ���  ���     �          �  #������?������������ ��������c��c�����    �  �  w������������  ;���  ����  ;���  ����  ;���  ���������c��c�����    �  �  w���������  �������  �  ����  �������  8  ������������c��c�����    �  �  w���������  �  8  ����������    �  �����������  � x� � �        ���  ���     �          �  #������?������������ ������������s��;���    �  �  w������������  ;���  ����  ;���  ����  ;���  �������������s��;���    �  �  w���������  �������  �  ����  �������  8  ����������������s��;���    �  �  w���������  �  8  ����������    �  �����������  c p � �        ���  ���     �          �  #������?������������ ������������{��{���    �  �  w������������  ;���  ����  ;���  ����  ;���  �������������{��{���    �  �  w���������  �������  �  ����  �������  8  ����������������{��{���    �  �  w���������  �  8  ����������    �  �����������  ! ` � �        ���  ���     �          �  #������?������������ �������������������    �  �  w������������  ;���  ����  ;���  ����  ;���  ��������������������    �  �  w���������  �������  �  ����  �������  8  �����������������������    �  �  w���������  �  8  ����������    �  �����������                   ���  ���     �          �  #������?������������ �������������������    �  �  w������������  ;���  ����  ;���  ����  ;���  ��������������������    �  �  w���������  �������  �  ����  �������  8  �����������������������    �  �  w���������  �  8  ����������    �  �����������                   ���  ���     �          �  #������?������������ �������������������    �  �  w������������  ;���  ����  ;���  ����  ;���  ��������������������    �  �  w���������  �������  �  ����  �������  8  �����������������������    �  �  w���������  �  8  ����������    �  �����������                   ���  ���     �          �  #������?������������ �������������������    �  �  w������������  ;���  ����  ;���  ����  ;���  ��������������������    �  �  w���������  �������  �  ����  �������  8  �����������������������    �  �  w���������  �  8  ����������    �  �����������                   ���  ���     �          �  #������?������������ ��           ��    �  �  w������������  ;���  ����  ;���  ����  ;���  ���           ��    �  �  w���������  �������  �  ����  �������  8  ������           ��    �  �  w���������  �  8  ����������    �  ����������� ���������������        ���  ���     �          �  #������?������������ ��               �����������������������������������������������������������������               �����������������������������������������������������������������               ���������������������������������������������������������������                  ����� ���?���������  ������������������������������������ ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                       �             @                                      ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������     � @       8   �  @pA      @              �  �$                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������     @ @      
 (   �   PA      @              
�  �
$                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������     U�wm�      
�#�� �  U�W]�     @              ������               ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ ������DUIT����  �"�� ����UTqU%���  �������������������*����������������� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      UDUIW       �"��    I�G]'                     ����                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      UEUIQ       �*��    UEQ$                     
�����$�                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ]Gui�       �;��    U�G]�                     ������                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                               ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                               ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ���             ������������������                                 ��       ����             ������������������                                 ��       ����             ������������������                                 ��       �  ��������������                  ���������������������������������� �������� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������               @                  �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@                  �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@                  �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@                  �                                        @ �����7�����������������������������޿�����������������������������������������������7�����������������������������޿�����������������������������������������������7�����������������������������޿������������������������������������������  �������������@   ` p (       �                                        @ �����������������������������������߿�����������������������������������������������������������������������������߿�����������������������������������������������������������������������������߿������������������������������������������  �������������@    � P         �                                        @ �����������������������������������ߧm��1���8�cN~3�q�c,nϗS���?������������������������������������������������ߧm��1���8�cN~3�q�c,nϗS���?������������������������������������������������ߧm��1���8�cN~3�q�c,nϗS���?�������������  �������������@ �����Gv�w      �                                        @ �����ձ�����k����������������������ߚ��]n����Z�]5��ٮ�}k���Mu���������������������ձ�����k����������������������ߚ��]n����Z�]5��ٮ�}k���Mu���������������������ձ�����k����������������������ߚ��]n����Z�]5��ٮ�}k���Mu����������������  �������������O�
���DET��T      �                                        @ �����5������o����������������������ߺ��A`���w��]v��۠��k�߷]}��������������������5������o����������������������ߺ��A`���w��]v��۠��k�߷]}��������������������5������o����������������������ߺ��A`���w��]v��۠��k�߷]}���������������  �������������@ :����ET��w      �                                        @ ������`�����o����������������������ߺ���_o����]w}�ۯ��k��]}����������������������`�����o����������������������ߺ���_o����]w}�ۯ��k��]}����������������������`�����o����������������������ߺ���_o����]w}�ۯ��k��]}����������������  �������������@ *���UT��A      �                                        @ ������o�����o����������������������޺��]n����Z�]u��ۮ��k���]u����������������������o�����o����������������������޺��]n����Z�]u��ۮ��k���]u����������������������o�����o����������������������޺��]n����Z�]u��ۮ��k���]u����������������  �������������@ 9J���wt�w      �                                        @ ������������������������������������n�cq���8�cv~7���lrϹ]���?�������������������������������������������������n�cq���8�cv~7���lrϹ]���?�������������������������������������������������n�cq���8�cv~7���lrϹ]���?�������������  �������������@                 �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@    0             �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@                  �                                        @ ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@                  �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �������������@                  �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������               @                  �                                        @ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��������������                  ���������������������������������� �������� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                  �C������ ������������ ���               ���������� ������������            /I�  �
�  ж?���-�;� ������������ /I�  �
�      �w� ������H�Q� ������������     ��w�             ���������� ������������     �              ���������� ������������     �                ���������� ������������     �              ���������� ������������     �              ���������� ������������     �              ���������� ���������������������          ���������� ����������������������          ���������� ����������������������          ���������� ����������������������          ?���������� ����������������������            ?���������� ����������������������      >      ����������������������@����������      ��     ������������          @                 x?�����?������������          @                 �         ��     ����� �����                                    ������������                    