�3{  �D d ��������������������������E��������������D�������C������H������������H��H���H��������H����������������������HC������������������������H�������B����������H������F��������H������H�����������H����������I����������H�����EI��������������C���H�����H���C���H�����B�����������������������������������������������II�������������������������G���I���������������������HD���GF�I���I��H�����CF�I���E�G��H��E��E�G�D��E��-��@
��
��@
l����@c����@�|
��@
e��w7
m��|@@1�*f��|@w����@�7
-�����������|
�7
l����?��@
w7
f��|@0�|
h�@1�|@0�@
m��|@7�o*
f�}6����@
��y@��@�������������|
4n��j.
gt@v�y@@��y*1�|@����@
u��@
r�~@m��?
d�@@���|@7
��?*r�|8�@��?*��@@��@*���@@@@���|���@
m������@��@*��@@��;m��?
�@��@*���|@��|@���>v�@|��|@7
��>7��{<5�@��>7��@@��@7��@@���@@m�|@m���|A@@@>��@7��@@
���@���>5�@��A7����@
��{@(���|7��@���@@
��{;��y@��@��|;��@@��@8��@@���@7(��@��|@7
��@8��@@m���?*(���|7��@��|;����|@��y@5����;
��@��@7��~@��>@��@@��@�������@;��@@��|@��?���@7
��@;���������A75����;
��@@��@��@��@��>@w�@��@��@��y@
���@��@@��|@@��@�������y<��������>@
��@��|@
(��y<���������|;w�@��@1�|@@��@��@��y@��@@��@��>*��@��y@�������@>���@��@@���@@��{@��������>?��?��A@4m����{@���@@��@��@��@��>*m��@��@@���@�@��@@�|@��|7��@��@�������?|�������@@��@@��|@	���@@@��|@��@��A@-����@��|@	��@@��@��@�|@��|;�������@@��~@��@��@@�A@��;���@��|���@���@��������@@��@@��}@��}@
m��@
(��@��|@0����@��}@��@@��@��@��>@��@�������@@��{@�@��@@�@;w�@��}@����3��}@��@��@@@��@@��@@���<��{@��|m��@���@@��?���?��@@��@�@��@;w�@��@@@��@@��>@����@@|@*�|@��{@m�����@��{@��@��y@�@@��@|����|��><	m��|��|@@��|
��|@���|��@|���@y���|@*�@��y@�@@��@;f���@@@@
b�@��>@j������><m�@��@;�@@�����������*
��@9m�����@@m��|
��@@������@������|@m��@@
b���@;�@@��@7���@@@7
7��@;
+x���@94�@@7*d@@����||���|@@@��@6j���|@7m�����|@7m��|@@����@�>;g|@7
7@@*d@@
7*m��@@
w�@7g�@6w@@


*;;*

7@7

8
*;;*
j���|@7

7@7

*7;�@7


@m�@@@*@@@@@@

@@@y
-���y
��y
��|
�����y
@@	&,m����?*5��@@m���@
1�����@@@5w���w*
5��q/
0clv����������������y7m�:
��@@����y*1m���j.
j���|@@
m�������@@m�����|
u�������������������;
1���?
��y@��@��;0��������=
t��@@7
m����|>@;7*m�������|
��������|@|�����|���@m���y*5��@;��@���@5���������|

��@@m��|@@7
���|@|���@
���~{>;96
,���@y���>����;���@*��@���?h��@@@@����?��@@��|@7
1��|@7
��|@��@@	$���@j��|7(�����@��|@�@���>6r��?m��@@��@@m�|@
f��@7
m��@��@@���@���<
4�����?*5��>@e�y@���{8��@��@@���|*
w�r�|@(��@@���|
��}@���@m�����>;���@@��@@��~<��|@��@@�����q*
@@w���0	��>@
��@@������j.

��|@5��>*������|@��@@�|@7���@��|?��?@������@@7*m����/
��>@��@@��������@
��y@
(��|;��||���@���y@���@���@��z@w�|@@���|A;7*3���|��|@��@@�������|@@��>@	���@��>>���?���@;���������?@��>@w��|@7��@@

m��@���@
��@@����|A;7*
��A<m��@���@@���?��|@*���������>@��@|���|@@7
��@@��@���@(��@@���}@
w�@;4��@���@7��@��@@���������{@��@��@@@7
��@@��@@��|@m��@@���{@m�@;��?��|@����@7m��@@@��~@���@���|��@@
w*
-��
m��?@���|m��|@@���>;	f�@7��@��>@
5���y@���y@���@��}@m���=
��@|��w*�@@���������|@7��������@@���@95�@75����@;m��@;���@;j��@��{@m����=�������@@�@@��������|@7
-������|@7w��@60�@6����@7g|@*��|@*�|@��A;m���@�������@@@@@j����|@7
j���|@7
g|@w@*m��|?*


77
b@@��@9
69<����|@@@*

*;@;*

*;;*



@m�@@

w@6	*;;*
@@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            