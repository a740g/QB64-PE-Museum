�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������{���������������������������������{���������������������������������{�������������������������������?������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������v�Ӈ��f?i����8{jS�ڔ�t�������v�Ӈ��f?i����8{jS�ڔ�t�������v�Ӈ��f?i����8{jS�ڔ�t�����?�����������������������������������~��Mw������]��{j��ڳ]u�k�������~��Mw������]��{j��ڳ]u�k�������~��Mw������]��{j��ڳ]u�k�����?�����������������������������������~��]w����.�A��z���]u��?������~��]w����.�A��z���]u��?������~��]w����.�A��z���]u��?����?�����������������������������������~��]w�wm����_���z���]u���������~��]w�wm����_���z���]u���������~��]w�wm����_���z���]u�������?�����������������������������������z��]w�u����]��}���v�]e��������z��]w�u����]��}���v�]e��������z��]w�u����]��}���v�]e������?������������������������������������{�]���v?.����8}�]�v�c����������{�]���v?.����8}�]�v�c����������{�]���v?.����8}�]�v�c�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������}����������������������������������}����������������������������������}��������������������������������?�����������������������������������}������������{���������������������}������������{���������������������}������������{�������������������?�����������������������������������9���������������������������������9���������������������������������9�������������������������������?�����������������������������������9�m�o�����v�ԧ���6����������9�m�o�����v�ԧ���6����������9�m�o�����v�ԧ���6��������?�����������������������������������U������u�꺿~��՚믶���]���������U������u�꺿~��՚믶���]���������U������u�꺿~��՚믶���]�������?�����������������������������������U������u���~��U�믶�s�]��������U������u���~��U�믶�s�]��������U������u���~��U�믶�s�]������?�����������������������������������mwk����u����~��U�믶���]���������mwk����u����~��U�믶���]���������mwk����u����~��U�믶���]�������?�����������������������������������mu�����u���z�����/����]���������mu�����u���z�����/����]���������mu�����u���z�����/����]�������?�����������������������������������}�n�k���_��{������7Wa��������}�n�k���_��{������7Wa��������}�n�k���_��{������7Wa������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������2��1������p��O�9���f?�������2��1������p��O�9���f?�������2��1������p��O�9���f?����?�����������������������������������tַ{~����]uu���}7��wַ]���������tַ{~����]uu���}7��wַ]���������tַ{~����]uu���}7��wַ]�������?�����������������������������������ְ{p�����u����w�v�]���������ְ{p�����u����w�v�]���������ְ{p�����u����w�v�]�������?�����������������������������������}ַ�n�����u}����w��uݷ����������}ַ�n�����u}����w��uݷ����������}ַ�n�����u}����w��uݷ��������?�����������������������������������uַ{n����]uu���]w��uַ]���������uַ{n����]uu���]w��uַ]���������uַ{n����]uu���]w��uַ]�������?������������������������������������ڸ�p���������w����?��������ڸ�p���������w����?��������ڸ�p���������w����?�����?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������'���a���q͸�����Ɵ�6����������'���a���q͸�����Ɵ�6����������'���a���q͸�����Ɵ�6����?�����������������������������������u��������u�����w]��}���ot�������u��������u�����w]��}���ot�������u��������u�����w]��}���ot�����?�����������������������������������u������u��������]�a����u�������u������u��������]�a����u�������u������u��������]�a����u�����?�����������������������������������u�������u�������w������u�������u�������u�������w������u�������u�������u�������w������u�����?�����������������������������������u�������u������]�]���u�?�����u�������u������]�]���u�?�����u�������u������]�]���u�?���?�������������������������������������������_a��������������������������_a��������������������������_a����������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?�����������������������������������>s1��|��bq�8�,i�?q��<����������>s1��|��bq�8�,i�?q��<����������>s1��|��bq�8�,i�?q��<��������?�����������������������������������u��n�۽��o����}k���鮳]}�[]�������u��n�۽��o����}k���鮳]}�[]�������u��n�۽��o����}k���鮳]}�[]�����?�����������������������������������t�7`�۽��-����k�����A}�[A�������t�7`�۽��-����k�����A}�[A�������t�7`�۽��-����k�����A}�[A�����?�����������������������������������u��o�۽��ۭ����k���뮷_}�[_�������u��o�۽��ۭ����k���뮷_}�[_�������u��o�۽��ۭ����k���뮷_}�[_�����?�����������������������������������u��n�۽��k����]k���뮷]}�[]�������u��n�۽��k����]k���뮷]}�[]�������u��n�۽��k����]k���뮷]}�[]�����?�����������������������������������>3���~��-��8�n����c}�[c������>3���~��-��8�n����c}�[c������>3���~��-��8�n����c}�[c����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������}���������������������������������}���������������������������������}�������������������������������?�����������������������������������}����������������������������������}����������������������������������}��������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������׍�i���������3=���S���������׍�i���������3=���S���������׍�i���������3=���S�������?������������������������������������u���V��]�������m��{�Mw��}j�������u���V��]�������m��{�Mw��}j�������u���V��]�������m��{�Mw��}j����?������������������������������������u��.�[��_�����v�m��{�]w��a��������u��.�[��_�����v�m��{�]w��a��������u��.�[��_�����v�m��{�]w��a�����?������������������������������������u����]��_u����mu���]w��]��������u����]��_u����mu���]w��]��������u����]��_u����mu���]w��]�����?������������������������������������u���V��]u�����mu�{-]w��]k������u���V��]u�����mu�{-]w��]k������u���V��]u�����mu�{-]w��]k���?������������������������������������_.�Y�������;=m���]���a��������_.�Y�������;=m���]���a��������_.�Y�������;=m���]���a�����?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������������������?���������������������������������?���������������������������������?�����������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?��������������������������������������������{��������������������������������{��������������������������������{���������������������?��������������������������������������������{��������������������������������{��������������������������������{���������������������?�������������������������������������M����8y�����'58{le������������M����8y�����'58{le������������M����8y�����'58{le��������?�����������������������������������u��5���o��{w�]����u��{k�w]��������u��5���o��{w�]����u��{k�w]��������u��5���o��{w�]����u��{k�w]������?�����������������������������������u��u���o��{w�A���t�z���]��������u��u���o��{w�A���t�z���]��������u��u���o��{w�A���t�z���]������?�����������������������������������u��u���ou�{w�_���u��z��w���������u��u���ou�{w�_���u��z��w���������u��u���ou�{w�_���u��z��w�������?�����������������������������������u��u϶�ou�{w�]���u��}ۭ�]��������u��u϶�ou�{w�]���u��}ۭ�]��������u��u϶�ou�{w�]���u��}ۭ�]������?�����������������������������������[�u߷o��}��c���5�}�m����������[�u߷o��}��c���5�}�m����������[�u߷o��}��c���5�}�m��������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������?����������������������������������?����������������������������������?����������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        