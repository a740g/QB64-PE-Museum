�3{  �D d ��������E����������������������E��������������������������������C������HD������HD�������C������C���F������H���HI������������������C��������������C����������������B���BB����������������������������II���IG��H�����������������E�����EI����I���������������H��������HB���I���I��������������HDC�������C���C��EC��EC���������B����������������������������������I��H����E��������B������I��I�������������E��������E�����I��I��H������������H������HHE��GG�GE��EE���EE���E�D�D��@
u|
u|
e�@
u|
4n��j.
4n��j.
5��q/
4n��j.
f��|@k�@
w7
o�@
w7
-�|
h�@@k�@
�����������������=
m�����|
4n��j.
5�������=
����@
��y*1�|@��y*1�|@0�@���@
r�@@4n��j.
��y*���@@�������@@����@���|���@
m������@
u��?@����@
�@��?@��;m��@
��;m��?
d�@@���|@��@|�������@
��;��@@�����?
m��@���@@m�|@m���|>@;7*���@
m��@*5�@��>?���@���>*(���@���>v�?@����@
��@����|>@;7*(���@��@@����}@��@���@7(��@��|@7
��}@��@;��?��|@����?*(���|74���?*(���|7��@@����|@��@��|@7
m���@*��@@����|@��@��|@��?���@7
��|@��@@��@@��@����>75����;s���>75����;
��@@��@��@�����@7
-�@
����A7��@@m��@��{@m��?��>@
��@��|@

��{@m��@@��|@@��@����|;w�@��@����|;w�@��@��@@��@��y@����|@
��@@����|;�������|���y@w��|��>?��?��A@5w��@��y@w��|@A���@��@��?��@��@��>@��@��@��@��>*��@@���@�?����>?5w��@7��@��@������|?��@���|@?y��|@��@��A@-�������@���|@@7�������@��@��@�|@��|@��@��@�|@��|7��@@��~@��@����>@-����@@��@��@���|>;7*��@��@@@
j��@
(��@��|@0����y}��?��@@@�������@��@��@��>@��@��@��@��A@��;��@@��{@�@����|@0����y@��@��@���~@
���@���|
��|m��@���@@��@{���@���|
m�@@@��@��@�@��@;w�@��@�@��@;w�@��@@��>@�������@@��@@��@�@���{@
��|@m��|
m��|��|@@��|
��|@A��|@m��|��y@�@��@y���|@*�@��@y���|@*�|@��@@��@;f���@��|
��|@@��@y�����><r�A@w�@m�����@@m��|
��@@��A@w�@��@;�@�|@m��@@
b��|@m��@@
b�@��@@��@7���@���|
��@@�k*
�|@m����@9f�?;
@@j���|@7m�����|@7��@<
777*d@�A;g|@7-�A;g|@7
7��@@
7*m��@@������|@7-�@@�A;g|��@61�@7
*;;*
j���|@7
d�@7
w@7

b@7

w�@@m�@@j���|@7

7�@7
@@*@@@@
@*@@@@@@@@@
@��|
�y
-���?��|
�y
�����m��>75�y@
%m�������>75�y*1������������=w=
w7
-������|
'���?@��@���������������?@��;4m���j.
j���|@��������@��|
w�@@��������@���|@7���@��������������|@7���@g��������=
t��@@7������������@
m�|@7��������@���@@
����@2�����|@@���@@
���@@����������|

��@@���@@@@��@��|@m��@@
���~{>?@@��@75��@,���@@��@75��@@���@@@@����?��@@��@@��@���@
m��|@7��@@���y@(��}@$���@���y@(��@@���@m��@@��@@��@?&w�|@@��|@��|@7
��@@���?;��{@
���@���@;��@@���@��@@���|��?����|@7m������@@
���|��@*��y?
��}@��@*��@@��}@��@@�����q�������|@
�����|?7�������@��y@��><
��|?��y@��@@��|?��?@��������������@
m���|@7
����������@@��@;��y@��@@��@@��{@w�|@@���|A;���|@@��@*)���@@
�������@��y@��@8��y@n�y@��@@��>@w��|@7��@@
��|@7��@;���@7����|>@@��@(��@6��@?f�@(��@@��@|���|@@7
��@@��@@��@;���@���}@j��@m��@+w�@<0��@m��@@��?��@@@7
��@@��@@m�|@*��|@���{@��|@��|@m�@9��|@��|@@���@���|��@@
��@|���@@
��y@	���>;	���&m��@@
f�?7���&m��@@��}@m���=
��@|����@���|@7m�A<���@95��������|@75�?7	5��������|@7t�{@m����=�����������|@7
e�@9���@6m������|@7
0�@6m������|@7
j�A<m���@����������|@7
0�?7	g|@j���|@7
w@*j���|@7
1�@9
69<����|m�|@7
w@6


*;;*

@
*;;*
w@6	*;;@@
@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            