��s  <
      PPPP��������������������          ����������������������������          pppp��������������������pppp          ����������������������������          ����������������������������          ����������������������������          pppp��������������������pppp          ����������������������������          ����                    ����          ����                ����@@@@          ����������������������������          ����������������������������          �����������ب���������������          �����������Ȩ���������������          pppp��������������������pppp          ����������������������������          pppp��������������������hhhh          ���������������𠠠���������          pppp��������pppp����pppp          ����                                  ������������������������pppp          ��������������������PPPP              �����������������������؈���          ��������PPPP    PPPP��������          ������������PPPP                      ����    @@@@@@@@����              ````                pppp          pppp����    @@@@����          pppp����0000����pppp          ����������������          ��������������������pppp          pppp��������������������pppp          ����                      pppp��������pppp��������pppp          pppp��������xxxx����pppp          pppp�������Ȩ�����������pppp                                                pppp��������������������pppp              PPPP����PPPP����PPPP              pppp��������pppp((((����pppp          ��������    @@@@XXXX����              PPPP����                          pppp����PPPP    XXXX����````              ����pppp����pppp����                  @@@@@@@@@@@@              @@@@        @@@@                      pppp                                  ����                              ����    ����                  pppp@@@@@@@@@@@@@@@@@@@@pppp          pppppppp          0000@@@@@@@@����@@@@@@@@0000          ````````          ����@@@@@@@@              PPPP����                              ````                                                      @@@@                                                    @@@@              ����@@@@        @@@@����          pppp����                          @@@@@@@@����                                                                        @@@@                                                                  