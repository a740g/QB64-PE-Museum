� {  �X \\]]^^_^_`__`aa   bbc         ffg   hihiijjjkkkklll   nno         rss   tuuvuvvvvwxwy     zz{{|||}}}}~~                       �����������       �����������     ���������������   ���������������   ���         ���     �����������     �������������     ���������������]]^^^___``aabbb   cdd         ghg   iijkkkkkllmmmmn   opp         sst   uvvwwwwwxxxxyz    {{|||}}}}~��                      �������������     �������������    ���������������   ���������������   ���         ���    �������������    ��������������    ���������������^__               dee         hhi         lmm         pqp         tuu   vww         zz{   |}|                                 ����       ����   ����       ����   ���                     ���         ���         ���   ����       ����   ���        ����   ���            __`               eff         iij         nnn         qqr         uvv   wwx          ||   ~~~                                 ���         ���   ���         ���   ���                     ���         ���         ���   ���         ���   ���         ���   ���            `aa               ffg         kjk         nnn         rrs         vvv   xyy          }|   ~~                                 ���         ���   ���         ���   ���                     ���         ���         ���   ���         ���   ���         ���   ���            aab               ggh         kll         oop         stt         wxx   yzz          }}   �                                 ���               ���         ���   ���                     ���         ���         ���   ���         ���   ���         ���   ���            bbc               hhi         lmm         pqq         ttu         xxy   {z{          ~   ���                                 ���               ���         ���   ���                     ���         ���         ���   ���         ���   ���         ���   ���            cdd               ijj         mmn         qrr         uuv         yzz   |||         ��   ���                                 ����              ���         ���   ���                     ���         ���         ���   ���         ���   ���        ����   ���            ddd               kjk         non         rrs         vvw         z{{   }|}~~}~���    ���                                  �������������    ���         ���   ����������              ���         ���         ���   ���         ���   ��������������    ���            eefffghhhih       kkl         oop         stt         xww         {||   ~}~~~������     ���������                             �������������   ���         ���   ����������              ���         ���         ���   ���������������   �������������     ���������      fgggghhhhii       llm         ppq         tuu         xxx         |}}   ~~~     ���       ���������                                      ����   ���         ���   ���                     ���         ���         ���   ���������������   ���     ���       ���������      ggh               mmn         qqr         vuv         yzy         }~~   ��     ���       ���                                             ���   ���         ���   ���                     ���         ���   ���   ���   ���         ���   ���     ���       ���            hii               noo         rrr         vww         {{{         ~~   ���      ���      ���                                             ���   ���         ���   ���                     ���         ���   ���   ���   ���         ���   ���      ���      ���            jii               opp         ttt         wxx         {{|         �   ���      ���      ���                                 ���         ���   ���         ���   ���                     ���         ���   ���   ���   ���         ���   ���      ���      ���            jjk               ppq         ttu         xxy         ||}         ���   ���      ���      ���                                 ���         ���   ���         ���   ���                     ���         ���   ���   ���   ���         ���   ���      ���      ���            kll               qrr         uuv         yyy         }~~         ���   ���       ���     ���                                 ���         ���   ���         ���   ���                     ���         ���   ���   ���   ���         ���   ���       ���     ���            llm               rrss       vvvw         zz{         ~       ����   ���       ���     ���                                 ����       ����   ����       ����   ���                     ���         ���� ����� ����   ���         ���   ���       ���     ���            nmn                tsttuuvvvvvww          {{|          ������������    ���       ���     ���������������                      �������������     �������������    ���                     ���          ������ ������    ���         ���   ���       ���     ���������������nno                 uuuuvwwwwwx           |}}           �����������     ���       ���     ���������������                       �����������       �����������     ���                     ���           ����   ����     ���         ���   ���       ���     ���������������                                                                                                                                                                                                 