�P  @                              0 0 @ 0 p 0   p p p  � � � ���  ���@���$� ;�?       ������������������������������������������������� � � � � � � � �����0�0�0�0�p�p�p�p��������                               �  0�0�0��`p���p�����D ?�{�?�0� ?�                           ��������������������������������?�?�?�?�            �����0�0�0�0������������������������                          @   ` `   p p p   p P p @ 8 x 8  < , <    >  � �  ���@���  ���������������������������������������������������������������������p�p�p�p�����0�0�0�0  �  ��� ��               
            	         ���@���  �p�p�p�p�p�p�p�p�����������������������������������������������������������������p�p�p�p�0�0�0�0          @���	 ��� ���   >  @ < | < @ 8 x 8   p p p  ` p ` @   ` `                   ���������0�0�0�0�����p�p�p�p������������������������������������������������������������                                  @���!�>��@@?��?�@p0xpp0 ` ``@ @ @                     ���������������������������������0�0�0�0� � � � � � � � ������������������������������������               �? ?� @���  ��� @���  � � �   p P p   p p p    0 0                  �����������������p�p�p�p�0�0�0�0��������� � � � ����������������������������������������                   � � � �   ���  ��� ���  ���� �  � � 	      �������������������������p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p��������