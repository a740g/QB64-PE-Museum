�P  (#� G �������������������������������������������������������������������������������������������������������������������������                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             ����������������������������� ����������������������������� �                           ������������������������������ �                            �                            �                           ��                            ����������������������������� ����������������������������� �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                         
 �                         
 �                         ������������������������������ �  8� �x� �        
 �  8� �x� �        
 �  8� �x� �        ������������������������������ �  �wp�>;�x;����   
 �  �wp�>;�x;����   
 �  �wp�>;�x;����   �������?��������������������� �  �}� >��?�8?�����  
 �  �|0 >�;�8?�����  
 �  �}� >��?�8?�����  �����c������_�������������� �  ��x?�~{����x��w���  
 �   `�8< |x��pxw �w���  
 �  ��x?�~{����x��w���  �����g���������������������� �  ��8~ ||����x��?�w���  
 �   a�8p x|���xp� 7�w���  
 �  ��8~ ||����x��?�w���  ������������������������|���� �   ��8� ||������ ?������  
 �   ��0� 8|������ ?p���8�  
 �   ��8� ||������ ?������  �����������������Ϝ������~?��� �  1��9��x|�������7��Ϲ�  
 �  1��1��x|����À����8  
 �  1��9��x|�������7��Ϲ�  ��������>�p �1��� �       $    @ 8 �� �  
 �                           
 �  0��q�y��9������?����|�  �����<?�?��  8~��p����� �    @�D   0 �  ��   
 �                           
 �  9��s��{��9���ǁ����<  �����<? ?��< 8|�������� �   @@   �     �  �  p   
 �                           
 �  9�����s��q���ǃ��w?�~  �����<> ?�8  8�?��������� �   @@`<   0 @@     0   
 �                           
 �  ?�������������?xw�?  �����|88 ?��0 8�?�� ������ �    ���C ` P@ @@$  
 �                           
 �  �����9�������?x�=�  �����|x ?�> `x�?��b����� �   ���|� �� @@0  
 �                           
 �  ������������?�>|���  �����|� ��~ px ������� �    <��  h�   
 �                           
 �  ��� ?�������<?���>  �����|�����#�|x���0G ���� �  �� q����8�<���   
 �                           
 �  �� ���s��;�|<ϸ��<  �����~�����~|��p������ �  ��� �� �c����8?�	�0  
 �                           
 �  ��� �� �c���8?�89�>  ���������������������������� �       �   c  p 8�<  
 �                           
 �       �   c  p 8�<  ������������������������������ �                   00   
 �                           
 �                   00   ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �     >  �        ��|     ������������������������������ �                           
 �                           
 �       �         �B     ������������������������������ �                           
 �                           
 �       �         �B     ������������������������������ �                           
 �                           
 �     p<�Hy��g���B     ������������������������������ �                           
 �                           
 �     �"�H�+ H� �|     ������������������������������ �                           
 �                           
 �     �"�H�� O���QB     ������������������������������ �                           
 �                           
 �     �"�H"�* H@�1B     ������������������������������ �                           
 �                           
 �     �"�0"�* H� �1B     ������������������������������ �                           
 �                           
 �     p<� y�$G��B     ������������������������������ �                           
 �                           
 �                        ������������������������������ �                           
 �                           
 �         � �              ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �     |        @   ���    ������������������������������ �                           
 �                           
 �     B        @   �     ������������������������������ �                           
 �                           
 �     B        @  "     ������������������������������ �                           
 �                           
 �     B�1����0H�A�
"     ������������������������������ �                           
 �                           
 �     |�J@IS(�QA""     ������������������������������ �                           
 �                           
 �     @�! �IR/�a�A"
"     ������������������������������ �                           
 �                           
 �     @��IR( QA""     ������������������������������ �                           
 �                           
 �     @�JAFR(�I�" �     ������������������������������ �                           
 �                           
 �     @�1��D�' D� ���     ������������������������������ �                           
 �                           
 �                         ������������������������������ �                           
 �                           
 �                         ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ��                            ����������������������������� ����������������������������� �                           ������������������������������ �                            �                            �                           ��                             ����������������������������� ����������������������������� �                           ��                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             �                             �                             ������������������������������                              ������������������������������                              ��������������������������������UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                  