�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ���� ��                        ���� ��                        ���� ��              ���������  ��@� 0                  ���� �� 0                  ���� �� 0                  ���� �� 0                        @�       0            ���� s��       0            ���� s��       0            ���� s��       0  ���������  ��@�       0            ���� y��       0            ���� y��       0            ���� y��       0               �  @�7�������;<��         ���� |��7�������;<��         ���� |��7�������;<��         ���� |��7�������;<�����������  ���@����6��l�ٳf�         ���� ~>����6��l�ٳf�         ���� ~>����6��l�ٳf�         ���� ~>����6��l�ٳf�            �� @���������3f��         ���� ~>���������3f��         ���� ~>���������3f��         ���� ~>���������3f�����������  ���@����3�����3f�`         ���� |�����3�����3f�`         ���� |�����3�����3f�`         ���� |�����3�����3f�`            �  @�0ٶ�6��l�ٳfͰ         ���� y��0ٶ�6��l�ٳfͰ         ���� y��0ٶ�6��l�ٳfͰ         ���� y��0ٶ�6��l�ٳfͿ���������  ��@�0ٶ�������<��         ���� s��0ٶ�������<��         ���� s��0ٶ�������<��         ���� s��0ٶ�������<��               @�                        ���� ��                        ���� ��                        ���� ��              ���������  ��@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������M����9��<�yN?�2Ɵ���D�1���������M����9��<�yN?�2Ɵ���D�1���������M����9��<�yN?�2Ɵ���D�1������?������������������������������������5m��ou֮�뽺�5��wֺou�M[}n���������5m��ou֮�뽺�5��wֺou�M[}n���������5m��ou֮�뽺�5��wֺou�M[}n������?������������������������������������um�}�t�����t���u�][a`���������um�}�t�����t���u�][a`���������um�}�t�����t���u�][a`������?������������������������������������umv}�u�������u��}ֺ�u�][]o���������umv}�u�������u��}ֺ�u�][]o���������umv}�u�������u��}ֺ�u�][]o������?�����������������������������������}umu�ou֮�뽺�u��uֺ�u�][]n��������}umu�ou֮�뽺�u��uֺ�u�][]n��������}umu�ou֮�뽺�u��uֺ�u�][]n������?�����������������������������������}um����9��=��v?����][a���������}um����9��=��v?����][a���������}um����9��=��v?����][a�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������0��������������������������������0��������������������������������0������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������p�q�>c=�����c��	�N�8�'1�������p�q�>c=�����c��	�N�8�'1�������p�q�>c=�����c��	�N�8�'1����?�����������������������������������k��鮺��}ֻ�{��j�u�������z�뮷�����k��鮺��}ֻ�{��j�u�������z�뮷�����k��鮺��}ֻ�{��j�u�������z�뮷���?������������������������������������.���~�}ۃ�{�a��u�녶���z���������.���~�}ۃ�{�a��u�녶���z���������.���~�}ۃ�{�a��u�녶���z������?������������������������������������������}ݿ�{W]��u��u�������������������}ݿ�{W]��u��u�������������������}ݿ�{W]��u��u����������?�����������������������������������k��뮺��}���{�]j�u��u����z�뮷�����k��뮺��}���{�]j�u��u����z�뮷�����k��뮺��}���{�]j�u��u����z�뮷���?������������������������������������p���>�~Y��|0����o����1�������p���>�~Y��|0����o����1�������p���>�~Y��|0����o����1����?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������q��������������������������������q��������������������������������q��������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������Sg�1�c������϶��÷�����������Sg�1�c������϶��÷�����������Sg�1�c������϶��÷�����?�����������������������������������u�뮺�v��[�n��m��|.�V�����ݷ�������u�뮺�v��[�n��m��|.�V�����ݷ�������u�뮺�v��[�n��m��|.�V�����ݷ�����?�����������������������������������u�믂�v��o�n��m���Y�ߪ��ݷ�������u�믂�v��o�n��m���Y�ߪ��ݷ�������u�믂�v��o�n��m���Y�ߪ��ݷ�����?�����������������������������������u�믾�v��w�n��m����Y�类�ݷ�������u�믾�v��w�n��m����Y�类�ݷ�������u�믾�v��w�n��m����Y�类�ݷ�����?�����������������������������������u��.��w>�[�n��m�{��V��ݮ����������u��.��w>�[�n��m�{��V��ݮ����������u��.��w>�[�n��m�{��V��ݮ��������?��������������������������������������]g�q��m��q����ݰ�������������]g�q��m��q����ݰ�������������]g�q��m��q����ݰ��������?������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������������������������?���������������������������������?���������������������������������?�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������?��������������������������������?��������������������������������?�����������������������������?�����������������������������������u��������������������������������u��������������������������������u������������������������������?�����������������������������������}��������������������������������}��������������������������������}������������������������������?�����������������������������������}����c�?�?41�~4�cm��2�c��������}����c�?�?41�~4�cm��2�c��������}����c�?�?41�~4�cm��2�c������?�����������������������������������>��V�]u��j�׮���Z�m���u�����������>��V�]u��j�׮���Z�m���u�����������>��V�]u��j�׮���Z�m���u���������?�����������������������������������u��0[�A���w`��Z�m��u�����������u��0[�A���w`��Z�m��u�����������u��0[�A���w`��Z�m��u���������?�����������������������������������u��7��_}��뿶��}�Z�m��uֺ���������u��7��_}��뿶��}�Z�m��uֺ���������u��7��_}��뿶��}�Z�m��uֺ�������?�����������������������������������u���V�]u���������Z�s��uֺ���������u���V�]u���������Z�s��uֺ���������u���V�]u���������Z�s��uֺ�������?������������������������������������>���c�7��?41�~7j�w���6�c���������>���c�7��?41�~7j�w���6�c���������>���c�7��?41�~7j�w���6�c������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?�������������������������������������q�8�|i�q�4�>�㇩��m��|f8��?�������q�8�|i�q�4�>�㇩��m��|f8��?�������q�8�|i�q�4�>�㇩��m��|f8��?���?�����������������������������������jk���Z������z��]w��Mm�m���[������jk���Z������z��]w��Mm�m���[������jk���Z������z��]w��Mm�m���[����?����������������������������������������n�.����{~��w��]m�m�|,o�����������n�.����{~��w��]m�m�|,o�����������n�.����{~��w��]m�m�|,o����?����������������������������������������v������{���w��]m�mu{��w�����������v������{���w��]m�mu{��w�����������v������{���w��]m�mu{��w����?�����������������������������������j���Z������z��]w��]s�mu{��[������j���Z������z��]w��]s�mu{��[������j���Z������z��]w��]s�mu{��[����?�������������������������������������q���|.���7{?,㇮��w�m�|.8g��������q���|.���7{?,㇮��w�m�|.8g��������q���|.���7{?,㇮��w�m�|.8g����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?��������������������������������������c=����|m�L6?��1��q���������������c=����|m�L6?��1��q���������������c=����|m�L6?��1��q����������?��������������������������������������]}m������������n�_���������������]}m������������n�_���������������]}m������������n�_����������?��������������������������������������A}m��y=��3�����`��/��������������A}m��y=��3�����`��/��������������A}m��y=��3�����`��/���������?�����������������������������������w��_}mu������u�����o�ۯ�����������w��_}mu������u�����o�ۯ�����������w��_}mu������u�����o�ۯ���������?�����������������������������������w��]}mu�����u�����n�[������������w��]}mu�����u�����n�[������������w��]}mu�����u�����n�[����������?��������������������������������������c}m�����m��6;��q��1��������������c}m�����m��6;��q��1��������������c}m�����m��6;��q��1���������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������?����������������������������������?����������������������������������?�������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������S���c�?��M���8�q�Ϙe1���������S���c�?��M���8�q�Ϙe1���������S���c�?��M���8�q�Ϙe1�������?�����������������������������������M���]}u�����5m���t�_��_k�n���������M���]}u�����5m���t�_��_k�n���������M���]}u�����5m���t�_��_k�n�������?�����������������������������������]���]a|���um���}�\/�_��`���������]���]a|���um���}�\/�_��`���������]���]a|���um���}�\/�_��`�������?�����������������������������������]����]}����umu��}�[���ۭo���������]����]}����umu��}�[���ۭo���������]����]}����umu��}�[���ۭo�������?�����������������������������������]���]]u����umu��u�[��_k�n���������]���]]u����umu��u�[��_k�n���������]���]]u����umu��u�[��_k�n�������?�����������������������������������]����a�?��um����\1�ߘm����������]����a�?��um����\1�ߘm����������]����a�?��um����\1�ߘm��������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        