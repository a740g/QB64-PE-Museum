�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������?�3��o&18��&o�>c�8��&18�������?�3��o&18��&o�>c�8��&18�������?�3��o&18��&o�>c�8��&18����?��������������������������������������w�����oo��j��ou����{�_o����������w�����oo��j��ou����{�_o����������w�����oo��j��ou����{�_o�����?����������������������������������������
�n����ou����{�n�����������
�n����ou����{�n�����������
�n����ou����{�n����?��������������������������������������}��w���m������ou�������m�����������}��w���m������ou�������m�����������}��w���m������ou�������m������?��������������������������������������u��w���m��j��u����z�_m����������u��w���m��j��u����z�_m����������u��w���m��j��u����z�_m�����?������������������������������������?����n�����?c����n��������?����n�����?c����n��������?����n�����?c����n�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������o����������������������������������o����������������������������������o����������������?���������������������������������������������������o����������������������������������o����������������������������������o����������������?�����������������������������������S�8���ӎ?p��s�)�ɌN?.Ɯq��������S�8���ӎ?p��s�)�ɌN?.Ɯq��������S�8���ӎ?p��s�)�ɌN?.Ɯq������?�����������������������������������M��{]u�Mu���[�of�������k���������M��{]u�Mu���[�of�������k���������M��{]u�Mu���[�of�������k�������?�����������������������������������]��}�u�]|��X7�n�ۅ�������������]��}�u�]|��X7�n�ۅ�������������]��}�u�]|��X7�n�ۅ�����������?�����������������������������������]����u��}���[��n��u��뵺����������]����u��}���[��n��u��뵺����������]����u��}���[��n��u��뵺��������?�����������������������������������]��{]u�]u���[�on��u��뻺���������]��{]u�]u���[�on��u��뻺���������]��{]u�]u���[�on��u��뻺�������?�����������������������������������]����Xݎ?���s���ۅ�?;��q��������]����Xݎ?���s���ۅ�?;��q��������]����Xݎ?���s���ۅ�?;��q������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������߱�������������������������������߱�������������������������������߱����������������?��������������������������������������������������.���������������������������������.���������������������������������.����������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������cO����c�����c�|8�46>���������cO����c�����c�|8�46>���������cO����c�����c�|8�46>������?�����������������������������������u��7���w��������mu��Z��ޛ�������u��7���w��������mu��Z��ޛ�������u��7���w��������mu��Z��ޛ�����?�����������������������������������u��w���������m��ou���������u��w���������m��ou���������u��w���������m��ou�������?�����������������������������������u��w��������u��m}�w�����������u��w��������u��m}�w�����������u��w��������u��m}�w���������?�����������������������������������u��w���w�����u��mu��Z��޻�������u��w���w�����u��mu��Z��޻�������u��w���w�����u��mu��Z��޻�����?�����������������������������������[cu�����������m�|8�46>��������[cu�����������m�|8�46>��������[cu�����������m�|8�46>������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������~��߫��}���������_�����������������~��߫��}���������_�����������������~��߫��}���������_��������?���������������������������������������������o{�������������������������������o{�������������������������������o{�������������������?�������������������������������������������{�o{�����������������������������{�o{�����������������������������{�o{�������������������?������������������������������������?��'^�}wo+�M��q��Ï��X��?��������?��'^�}wo+�M��q��Ï��X��?��������?��'^�}wo+�M��q��Ï��X��?�����?�������������������������������������vj��^����j��5oi����w���WM���������vj��^����j��5oi����w���WM���������vj��^����j��5oi����w���WM�����?�������������������������������������v�����woj�u����������]���������v�����woj�u����������]���������v�����woj�u����������]�����?�����������������������������������u������;�oj��u�ۮ���������������u������;�oj��u�ۮ���������������u������;�oj��u�ۮ�������������?�����������������������������������u�����~���oj��uok����w���W]�������u�����~���oj��uok����w���W]�������u�����~���oj��uok����w���W]�����?����������������������������������������^����k�u�����Ï�V��ݿ������������^����k�u�����Ï�V��ݿ������������^����k�u�����Ï�V��ݿ�����?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������������n��������������������������������n��������������������������������n������������?�����������������������������������1�v��D�1�㌱��6?������c���������1�v��D�1�㌱��6?������c���������1�v��D�1�㌱��6?������c�������?�����������������������������������n���M[}n��u��ݵ���}���������������n���M[}n��u��ݵ���}���������������n���M[}n��u��ݵ���}�������������?�����������������������������������n���][a`��}��ߵ��z���������������n���][a`��}��ߵ��z���������������n���][a`��}��ߵ��z�������������?�����������������������������������n���][]o��}��ߵ���wn�������������n���][]o��}��ߵ���wn�������������n���][]o��}��ߵ���wn�����������?�����������������������������������n���][]n��u������ﯮ��������������n���][]n��u������ﯮ��������������n���][]n��u������ﯮ������������?�����������������������������������q���][a��Ꮁ���67�����������������q���][a��Ꮁ���67�����������������q���][a��Ꮁ���67���������������?������������������������������������������������������������������������������������������������������������������������������������������?��������������������������������������������������?����������������������������������?����������������������������������?�����������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������>��_}������_���������������������>��_}������_���������������������>��_}������_�������������������?�����������������������������������u����{����������������������������u����{����������������������������u����{��������������������������?�����������������������������������u�{��{���������ݿ�����������������u�{��{���������ݿ�����������������u�{��{���������ݿ���������������?�����������������������������������u�{��y��l=�8T��ݧ~0�MN��������u�{��y��l=�8T��ݧ~0�MN��������u�{��y��l=�8T��ݧ~0�MN������?�����������������������������������;���{u�뫽w�S]�ݚ��]55�����������;���{u�뫽w�S]�ݚ��]55�����������;���{u�뫽w�S]�ݚ��]55���������?�����������������������������������w۽w�{u���vW]�����Auu�����������w۽w�{u���vW]�����Auu�����������w۽w�{u���vW]�����Auu���������?�����������������������������������w�=w�{u�뫽u�W]������_uu���v�������w�=w�{u�뫽u�W]������_uu���v�������w�=w�{u�뫽u�W]������_uu���v�����?�����������������������������������u����{u�뫽u�W]�w���]uu���w������u����{u�뫽u�W]�w���]uu���w������u����{u�뫽u�W]�w���]uu���w����?�����������������������������������7��x{��l=�Waw��0�uv�������7��x{��l=�Waw��0�uv�������7��x{��l=�Waw��0�uv�����?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������������������?����������������������������������?����������������������������������?��������?������������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������������}������������_�������������������}������������_�������������������}������������_������?�����������������������������������������������}w�����������_��������������������}w�����������_��������������������}w�����������_������?����������������������������������������������׻w�����������_�������������������׻w�����������_�������������������׻w�����������_������?�����������������������������������S��~6�ӛ��w���p��1��X�[�������S��~6�ӛ��w���p��1��X�[�������S��~6�ӛ��w���p��1��X�[�����?�����������������������������������Mw�k�ַMj鿻������]n���}[�������Mw�k�ַMj鿻������]n���}[�������Mw�k�ַMj鿻������]n���}[�����?�����������������������������������]w��<�]�뿻�w���.�]n����[�������]w��<�]�뿻�w���.�]n����[�������]w��<�]�뿻�w���.�]n����[�����?�����������������������������������]w�������뿃�w�����]n����[�������]w�������뿃�w�����]n����[�������]w�������뿃�w�����]n����[�����?�����������������������������������]w��ַ]j�}}w����Yn���]\��������]w��ַ]j�}}w����Yn���]\��������]w��ַ]j�}}w����Yn���]\������?�����������������������������������]���~6�ݛ�}}���p�e���X�]��������]���~6�ݛ�}}���p�e���X�]��������]���~6�ݛ�}}���p�e���X�]������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        