�P  X  �  ���  ���  ���  ��    8  888x  8x8x88  88888x  8x8x8p  8p8p80  80809�  9�9�                                          �   � ��  ���  ���  ���  ���  ���  ��                    �  ��                                            �   � ��  ��8  88<  <<8  888  880  00 `   ` ` `   ` ` �   � ��  ��     �  ��?�  ?�?�                                     �   � ��  ���  ��<  <<8  88 x   x x 0   0 0 �   � ��  ���  ��x  xx <   < < x   x x�  ��                                  