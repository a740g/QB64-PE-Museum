�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������?����?���������������������������?����?���������������������������?����?�����������������������?���?����?������������������������?��������?�������������������������?��������?�������������������������?��������?�����������������������?�?��������?���������������������������������?����������������������������������?����������������������������������?�����������������������?����������?���������������������������0�����1����������������������������0�����1����������������������������0�����1�����������������������?����0�����1������������������������fL�>I��̙$�������������������������fL�>I��̙$�������������������������fL�>I��̙$�����������������������?�fL�>I��̙$������������������������&@�0I��̙3�������������������������&@�0I��̙3�������������������������&@�0I��̙3�����������������������?�&@�0I��̙3������������������������&O�&I��̙9�������������������������&O�&I��̙9�������������������������&O�&I��̙9�����������������������?�&O�&I��̙9������������������������&L�&I��̙$�������������������������&L�&I��̙$�������������������������&L�&I��̙$�����������������������?�&L�&I��̙$������������������������`��0L����1�������������������������`��0L����1�������������������������`��0L����1�����������������������?�`��0L����1�������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������o���������������������������������o���������������������������������o�������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������)��ߍ;[S����le��>c�lm�C�q��������)��ߍ;[S����le��>c�lm�C�q��������)��ߍ;[S����le��>c�lm�C�q�����?�����������������������������������k��꺿��[Mu��{k��w������]���������k��꺿��[Mu��{k��w������]���������k��꺿��[Mu��{k��w������]�������?������������������������������������������U]��z��������]�������������U]��z��������]�������������U]��z��������]����?�����������������������������������������u�U]}��z��~�}������]������������u�U]}��z��~�}������]������������u�U]}��z��~�}������]����?����������������������������������������u���u��}ۭ��u������]��������������u���u��}ۭ��u������]��������������u���u��}ۭ��u������]�������?������������������������������������.�����ݍ��}�m��c�ln�C�q��������.�����ݍ��}�m��c�ln�C�q��������.�����ݍ��}�m��c�ln�C�q�����?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������������������x?����_���������������������������x?����_���������������������������x?����_�����?����  ������������������������������������������������{���������������������������������{���������������������������������{�����������?����  ������������������������������������������������{���������������������������������{���������������������������������{�����������?����  ����������������������������������xᅎ|8�lq��o�8xm�q_�������������xᅎ|8�lq��o�8xm�q_�������������xᅎ|8�lq��o�8xm�q_�����?����  ��������������������������������=��w]uu��[k���o��{��j������������=��w]uu��[k���o��{��j������������=��w]uu��[k���o��{��j������?���� <��������������������������������=��w]u��Z� ��������������������=��w]u��Z� ��������������������=��w]u��Z� ��������������?����<��������������������������������=��w]u}�ګ���u����������������=��w]u}�ګ���u����������������=��w]u}�ګ���u����������?����<��������������������������������=��w]uu��]ۮ��ou�{���������������=��w]uu��]ۮ��ou�{���������������=��w]uu��]ۮ��ou�{���������?����
<��������������������������������=��xᅎ|8��q��o��|m���������������=��xᅎ|8��q��o��|m���������������=��xᅎ|8��q��o��|m���������?����<�����������������������������������������������������������������������������������������������������������������������������������?���� <��������������������������������}���������������������������������}���������������������������������}���������������������������?���� <�����������������������������������������������������������������������������������������������������������������������������������?����������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������8�~3�q�c���=�2�p���������������8�~3�q�c���=�2�p���������������8�~3�q�c���=�2�p�������?����  ������������������������������������Z��ٮ��mw��k��ֻ��M���������������Z��ٮ��mw��k��ֻ��M���������������Z��ٮ��mw��k��ֻ��M�����?����  ������������������������������������Z��۠��m�
�U�x.�]���������������Z��۠��m�
�U�x.�]���������������Z��۠��m�
�U�x.�]�����?����  ������������������������������������Z��ۯ��m���Uֻ��]���������������Z��ۯ��m���Uֻ��]���������������Z��ۯ��m���Uֻ��]�����?����  ������������������������������������Z��ۮ��mw�����ۮ�]���������������Z��ۮ��mw�����ۮ�]���������������Z��ۮ��mw�����ۮ�]�����?����  �������������������������������  �8k�7���m���>�6�p�����������  �8k�7���m���>�6�p�����������  �8k�7���m���>�6�p������?������������������������������������������������������������������������������������������������������������������������������������������?����  ��������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?����  ��������������������������������������������������������������������������������������������������������������������������������?����  �������������������������������������ߍ;|q����q�N8c������������������ߍ;|q����q�N8c������������������ߍ;|q����q�N8c�������?����  ����������������������������������������{����ٮ���]�����������������������{����ٮ���]�����������������������{����ٮ���]���������?����  ���������������������������������������{�۠��A��������������������{�۠��A��������������������{�۠��A�������?����  ��������������������������������������u�{�ۯ���_��u�����������������u�{�ۯ���_��u�����������������u�{�ۯ���_��u�����?����  �������������������������������������u������ۮ���]��u����������������u������ۮ���]��u����������������u������ۮ���]��u�����?����"���������������������������������������q������c��������������������q������c��������������������q������c�������?�������������������������������������*���������������������������������*���������������������������������*���������������������������?����"���������������������������������o����������������������������������o����������������������������������o���������������������������?���� ���������������������������������o����������������������������������o����������������������������������o���������������������������?���� �������������������������������A��������������������������������A��������������������������������A���������������������������?����@���������������������������������������������������������������������������������������������������������������������������?���� ���������������������������������������������������������������������������������������������������������������������������?���� ����������������������������������o�Nf4�~3��N4Ꮨ�q�㍌�������������o�Nf4�~3��N4Ꮨ�q�㍌�������������o�Nf4�~3��N4Ꮨ�q�㍌������?���� �����������������������������������5��]u����7�]w�{���uu���������������5��]u����7�]w�{���uu���������������5��]u����7�]w�{���uu������?����  �����������������������������������v�_����v]�{���uu���������������v�_����v]�{���uu���������������v�_����v]�{���uu������?����  �����������������������������������wm�_}���u�]�{���uu���������������wm�_}���u�]�{���uu���������������wm�_}���u�]�{���uu������?����  �����������������������������������u��]u����u�]w�{���uu���������������u��]u����u�]w�{���uu���������������u��]u����u�]w�{���uu������?����  �����������������������������������vvc�~7��va���q�㍍���������������vvc�~7��va���q�㍍���������������vvc�~7��va���q�㍍������?����  �������������������������������  ��������������������������������  ��������������������������������  ���������������������������?������������������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������������?����  �����������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        