�P�pI� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                               ��                               ��                               ��                               ��                               ��                               ��                               ��              ����������������@����                         �����                         �����                         �����                         @��`                         s���`                         s���`                         s���`        ����������������@��                          y���                          y���                          y���                          @����8                       |�����8                       |�����8                       |�����8      ����������������@����6l                       ~>����6l                       ~>����6l                       ~>����6l                       @���60                       ~>���60                       ~>���60                       ~>���60      ����������������@���6                       |����6                       |����6                       |����6                       @��l�6l                       y���l�6l                       y���l�6l                       y���l�6l      ����������������@�ϳǙ�8                       s��ϳǙ�8                       s��ϳǙ�8                       s��ϳǙ�8                       @�                               ��                               ��                               ��              ����������������@�                               ��                               ��                               ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������                                 �޿�������������������������������޿�������������������������������޿�������������������������������                                 �߿�������������������������������߿�������������������������������߿�������������������������������                                 �߬m��c<��?������������������������߬m��c<��?������������������������߬m��c<��?������������������������                                 �߫��]]}��u������������������������߫��]]}��u������������������������߫��]]}��u������������������������                                 �߫���]}��u������������������������߫���]}��u������������������������߫���]}��u������������������������                                 �߫���]}��u������������������������߫���]}��u������������������������߫���]}��u������������������������                                 �ޫ��]]}��u������������������������ޫ��]]}��u������������������������ޫ��]]}��u������������������������                                 ��n��c~�ㅿ�������������������������n��c~�ㅿ�������������������������n��c~�ㅿ������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��    |    �    |    �    |    ���    |    �    |    �    |    ���    |    �    |    �    |    ��?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    �������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    �������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    �������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    �������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    �������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    �������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������     B         B         B    ����������������������������������������������������������������������������������������������������������?����������?����������?��������������������������������������������������������������������������������������������������������������������                                 ��    |    �    |    �    |    ���    |    �    |    �    |    ���    |    �    |    �    |    ��?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?�����������������    ������    ������    ���    }�����������    �    }��������    |    �    }������������������?����������?����������?��������������������������������������������������������������������������������������������������������������������?����������?����������?��������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������     �����������������������������     �����������������������������     ��                          ���������������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ����                   ?���������������                   ?����     �����                   ?����     ��  ��������������������        ����                   ?���������������                   ?����     �����                   ?����     ��  @                            ���������������������������������������������������������������     �����������������������������     ��  ��������������������        ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ����                   ?���������������                   ?����     �����                   ?����     ��  ��������������������        ����                   ?���������������                   ?����     �����                   ?����     ��  @                            ���������������������������������������������������������������     �����������������������������     ��  ��������������������        ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ����                   ?���������������                   ?����     �����                   ?����     ��  ��������������������        ����                   ?���������������                   ?����     �����                   ?����     ��  @                            ���������������������������������������������������������������     �����������������������������     ��  ��������������������        ���������������������������������������������������������������     �����������������������������     ��                               ���������������������������������������������������������������     �����������������������������     ��                               ����������������������������������������������������������������������������������������������������������                          ����������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������          �����������������������          �����������������������          ��                                 ����������������������������������������������������������������������������������������������������������                    ����������������������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     �����_�������������������������������_�������������������������������_���������������������������                         !     ��������������������������z������������������������������z������������������������������z�����                         !     ��������������������������z������������������������������z������������������������������z�����                         !     ���]��Xc3�5����1��0����N8����z������]��Xc3�5����1��0����N8����z������]��Xc3�5����1��0����N8����z����                         !     ���]k�W]m��u~��n�]u�_���5�_���z������]k�W]m��u~��n�]u�_���5�_���z������]k�W]m��u~��n�]u�_���5�_���z����                         !     ���]��WAw��|��n�_|_���u�_���z�������]��WAw��|��n�_|_���u�_���z�������]��WAw��|��n�_|_���u�_���z�����                         !     ���]��W_{��}~��n�_}�_���u�����z�������]��W_{��}~��n�_}�_���u�����z�������]��W_{��}~��n�_}�_���u�����z�����                         !     ��]Yk�W]m��u���n�]u�_��]u�_���z������]Yk�W]m��u���n�]u�_��]u�_���z������]Yk�W]m��u���n�]u�_��]u�_���z�����                         !     ��ae��Xcs�5����c�0����v8�����������ae��Xcs�5����c�0����v8�����������ae��Xcs�5����c�0����v8����������                         !     ����������������������������������������������������������������������������������������������������                         !     �������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������������������������������������������������������������������������������������������                         !     ����������������������          �����������������������          �����������������������          ��                    ����������������������������������          �����������������������          �����������������������          ��                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                         	 ��������������������������������������������������      ��                                                                                                                             	 ������  ������  ������        ��        ��������������  ������  ������                                                                                                                              