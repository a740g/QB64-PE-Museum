�P  �> P -                                              �         �         �         �         �         �         �         �         �         �         �                   �         �        �                   �         �        ;�                   �         �       �                   �         �       ��                   �         �       ��                   �         �       ��                   �         �       ��                   �         �       ��                   �         �       Ā                   �         �       ��                   �         �        �                   �         �         �                   �         �         �                   �         �         �                                               �����               �����     �����                         �����     �����                         �����     �����              �����    �����                        �����    �����               ����     �����    �����               ����     �����    �����                        �����    �����              wwww     �����    �����              wwww@    �����    �����              wwww`    �����    �����              wwwwp    ?�����    ?�����              wwwwp    �����    �����              7wwwwt    ������    ������              tp@   �������  �������   ���    tp@   �������  ����   @   tp@   �������  ����   @   tp@@  �������  ����   @   tp@`  �������  ����   @   tp@p  ?�������  ?�������   ���   tp@p  �������  ����   @   7tp@t  ��������  �����   @   wtp@v ���������������  @            ���������������  @  ������������������������  ���  ������������������������                                          �����        �����                     ]����       �����       �����                     �����       �����       �����                    �����       �����       �P - �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������� �������� �������� �������� �������� �������� �������� �������� �������� �������� �������� �������� �������� �������� �������� ����������������������������������������;��������;��������;��������;���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������UUUU�����UUUU�����UUUU�����UUUU�����UUUU�����UUUU�����UUUU�����UUUU�����    �����    �����    �����    �����UUUU�����UUUU�����UUUU�����UUUU�����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    ?�����    ?�����    ?�����    ?�����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    ����      ����      ����      ����      ����      ���      ���      ���      ���      ?���      ?���      ?���      ?���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ��        ��        ��        ��        ��        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �~��?���  ?����������  ?�~��?���               >0f��3`��  ?����������  ?�~��?���               ?�~��?���  ?����������  ?�~��?���               >0f��3`��  ?����������  ?�~��?���    P                               ������������������������������������          ���������������������������          ���������������������������          ���������������������������                                                  x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?�������?����          x���������?�������?����          ��?���������������?�����          x��3�`������������?�����          ��?���������������?�����          x��3�`������������?�����          ���������������������������          x��3�`������������?�����          ��?���������������?�����          x��3�`������������?�����          ��?���������������?�����          x��3�`������������?�����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          ������������������?����          x����������������?����          ���������?�������������          x���`����?�������������          ���������?�������������          x���`����?�������������          ���������������������������          x���`����?�������������          ���������?�������������          x���`����?�������������          ���������?�������������          x���`����?�������������          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x�������������������������          �����������?������?����          x���������?������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���������������������������          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ��?���������������?����          x��3`�������������?����          ���x����x����x� ��?��� x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          x        ������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����