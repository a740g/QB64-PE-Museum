�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������_������������������������������_������������������������������_������?������������������������������������������w�������o���������������������w�������o���������������������w�������o������������?������������������������������������������w�������o���������������������w�������o���������������������w�������o������������?�����������������������������������|�'�c�3�w��N?p��)�����8WX]�������|�'�c�3�w��N?p��)�����8WX]�������|�'�c�3�w��N?p��)�����8WX]�����?��������������������������������������]mt�ݏ�{5���_f�ڻ���WW]����������]mt�ݏ�{5���_f�ڻ���WW]����������]mt�ݏ�{5���_f�ڻ���WW]�����?�����������������������������������}���Am��w�{t��_n�ڃ���Z�]�������}���Am��w�{t��_n�ڃ���Z�]�������}���Am��w�{t��_n�ڃ���Z�]�����?�����������������������������������}���_m}��w�{u����_n�ڿ���Z�]u������}���_m}��w�{u����_n�ڿ���Z�]u������}���_m}��w�{u����_n�ڿ���Z�]u����?�����������������������������������}���]mu��w�{u���_n�ڻ���]�Yu������}���]mu��w�{u���_n�ڻ���]�Yu������}���]mu��w�{u���_n�ڻ���]�Yu����?�����������������������������������}���cm�����v?��߮������]�e�������}���cm�����v?��߮������]�e�������}���cm�����v?��߮������]�e�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������������.��������������������������������.��������������������������������.�������������������?������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������&18�����X���S1��3ɌN?��������&18�����X���S1��3ɌN?��������&18�����X���S1��3ɌN?������?�����������������������������������o��zku���M�����Mn��ou����߆��������o��zku���M�����Mn��ou����߆��������o��zku���M�����Mn��ou����߆������?�����������������������������������n�z�u���]���]`��tۅ����������n�z�u���]���]`��tۅ����������n�z�u���]���]`��tۅ��������?�����������������������������������m����u���]��]o���u��u�����������m����u���]��]o���u��u�����������m����u���]��]o���u��u���������?�����������������������������������m��z�u���]��]n��ou��u�߾��������m��z�u���]��]n��ou��u�߾��������m��z�u���]��]n��ou��u�߾������?�����������������������������������n��덶�X��߱�]���7ۅ�7��������n��덶�X��߱�]���7ۅ�7��������n��덶�X��߱�]���7ۅ�7������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������A���x7����������������������������A���x7����������������������������A���x7������������������?��������������������������������������������v��{׻���������������������������v��{׻���������������������������v��{׻����������������?���������������������������������������������v��{׻����������������������������v��{׻����������������������������v��{׻����������������?������������������������������������������1��v��{׻�|�g�������������������1��v��{׻�|�g�������������������1��v��{׻�|�g����������?�����������������������������������u������~�ݎ��x7��k�����k�����������u������~�ݎ��x7��k�����k�����������u������~�ݎ��x7��k�����k���������?�����������������������������������p�����p��v�U{����=��h?����������p�����p��v�U{����=��h?����������p�����p��v�U{����=��h?��������?�����������������������������������~n����n��v�U{������o��k�����������~n����n��v�U{������o��k�����������~n����n��v�U{������o��k���������?�����������������������������������u������n��v��{���뽭���k�����������u������n��v��{���뽭���k�����������u������n��v��{���뽭���k���������?����������������������������������������{�p����{�{��}�w�lw���������������{�p����{�{��}�w�lw���������������{�p����{�{��}�w�lw��������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������o��������������������������������o��������������������������������o�������������������������?��������������������������������������غ뷷������������������������������غ뷷������������������������������غ뷷�������������������������?��������������������������������������޾ﷷ������������������������������޾ﷷ������������������������������޾ﷷ�������������������������?������������������������������������&;^�﷔��8Ӈ���8���&蟌����������&;^�﷔��8Ӈ���8���&蟌����������&;^�﷔��8Ӈ���8���&蟌�������?������������������������������������o�^�w�]�u�Mw�[���{jj��o��m��������o�^�w�]�u�Mw�[���{jj��o��m��������o�^�w�]�u�Mw�[���{jj��o��m�����?������������������������������������n^�ﷷA��]w�[���{j���o��m��������n^�ﷷA��]w�[���{j���o��m��������n^�ﷷA��]w�[���{j���o��m�����?������������������������������������m�^�ﷷ_�}�]w������j���ou�m��������m�^�ﷷ_�}�]w������j���ou�m��������m�^�ﷷ_�}�]w������j���ou�m�����?�����������������������������������}m�޺뷷]�u�]w�[���{j���ou�s�������}m�޺뷷]�u�]w�[���{j���ou�s�������}m�޺뷷]�u�]w�[���{j���ou�s�����?�����������������������������������}n��w�c�8݆��o���j��+o��w�������}n��w�c�8݆��o���j��+o��w�������}n��w�c�8݆��o���j��+o��w�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������~�����������q�?�������������������~�����������q�?�������������������~�����������q�?����?������������������������������������������������������������뮏��������������������������������뮏��������������������������������뮏�����?���������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������q����Ϗ������cN8�?�����������q����Ϗ������cN8�?�����������q����Ϗ������cN8�?�������?�����������������������������������k�y���[뷷_��}�[]�u�]5�z��}��������k�y���[뷷_��}�[]�u�]5�z��}��������k�y���[뷷_��}�[]�u�]5�z��}������?�������������������������������������{�����_�뽸[A��Au�{������������{�����_�뽸[A��Au�{������������{�����_�뽸[A��Au�{��������?������������������������������������w�����뷷_w뽷[_�}�_u���{����������w�����뷷_w뽷[_�}�_u���{����������w�����뷷_w뽷[_�}�_u���{�������?�����������������������������������j�{���Z�Ϸ_w뽷[]�u�]u�z�����������j�{���Z�Ϸ_w뽷[]�u�]u�z�����������j�{���Z�Ϸ_w뽷[]�u�]u�z���������?����������������������������������������߸߇�}�[c�cv8�>`�������������߸߇�}�[c�cv8�>`�������������߸߇�}�[c�cv8�>`������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������?����������������������������������?����������������������������������?������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������?��?���������0����������������?��?���������0����������������?��?���������0����?�������������������������������������������_��������������u����������������_��������������u����������������_��������������u������?�������������������������������������������߷������������������������������߷������������������������������߷��������������������?�����������������������������������~2&��Ɏ��w��߿�߿߿|�'����������~2&��Ɏ��w��߿�߿߿|�'����������~2&��Ɏ��w��߿�߿߿|�'��������?����������������������������������������������>?��?�߿����7�����������������>?��?�߿����7�����������������>?��?�߿����7����?�����������������������������������}����ۆ�]����m��}����w�������}����ۆ�]����m��}����w�������}����ۆ�]����m��}����w�����?�����������������������������������}������v�[��=߿߿߿}�����w�������}������v�[��=߿߿߿}�����w�������}������v�[��=߿߿߿}�����w�����?�����������������������������������}�����[w7W���߿�߿߿}����u�������}�����[w7W���߿�߿߿}����u�������}�����[w7W���߿�߿߿}����u�����?�����������������������������������~6�+�[�x��?��?���}�����8�������~6�+�[�x��?��?���}�����8�������~6�+�[�x��?��?���}�����8�����?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        