�  X           <<< fff fff fff fff fff fff fff <<<                        xxx                              <<< fff     000 ``` ~~~                       <<< fff      fff <<<                          <<< <<< lll ~~~                         ~~~ ``` ``` ||| fff   fff <<<                       <<< fff ``` ``` ||| fff fff fff <<<                       ~~~      000 000 000                       <<< fff fff fff <<< fff fff fff <<<                       <<< fff fff fff >>>   fff <<<            