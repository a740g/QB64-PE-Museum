�P   N � ���������������������������������������������������������������������������������������������������������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �?������������������������������?����������������������������� ��                            ������������������������������� �                             �                              ��                            ��                             �/������������������������������/����������������������������� ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                        ����(�(                        ����( ��                        ���������������������������������� �(                        ����(�(                        ����( ��                        �������������������������������?�� �( �9��O>�Bp              ����(�( �9��O>�Bp              ����( �� �9��O>�Bp              ��?���������������������������� �� �( �DD(P��b�              ����(�( �DD(P��b�              ����( �� �DD(P��b�              � ���������������������������� �� �( �@D(P�b�              ����(�( �@D(P�b�              ����( �� �@D(P�b�              � ���������������������������� �� �( �@D(P�R�              ����(�( �@D(P�R�              ����( �� �@D(P�R�              � ���������������������������� �� �(                        �� (�(                        �� ( �� �8G�P�Rp              � ���������������������������� �� �(                        �� (�(                        �� ( �� �D(P�J              � ���������������������������� �� �(                        �� (�(                        �� ( �� �D(P�F              � ���������������������������� �� �(                        �� (�(                        �� ( �� �DD(P��F�              � �����������������������������?�� �(                          � (�(                          � ( �� �8D'��Bp              ��?������������������������������� �(                          � (�(                          � ( ��                        ���������������������������������� �(                            (�(                            ( ��                        ����������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ����������������������������� �(                            (�(                            ( �� �              � P    ��������������������������� �(                            (�(                            ( �� "    �	       � � �   ��������������������������� �(                            (�(                            ( �� "    �	       � � �   ����8�0��?�bq�?1�q�N?)����� �(                            (�(                            ( �� "��'��c��������f   �����}�W]~��k�ﭮ��n���5�kk���� �(                            (�(                            ( �� #(�(���	�ARQ �Q� ��   �����}�P_~���>�-��n���tk����� �(                            (�(                            ( �� "/�(���	��_��_���D   �������W�~����뭯��n���u�k����� �(                            (�(                            ( �� "((� �	RP@�P� �$   �����}�W]~���뭮��n���u�kk���� �(                            (�(                            ( �� "(�(���	ARQ �Q� ��   ������0����-��?��q�v?k����� �(                            (�(                            ( �� "'�'@����N�N����b   ������������������������������� �(                            (�(                            ( ��                           ������������������������������ �(                            (�(                            ( ��           �               ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( ��        �       �A      ������������������������������� �(                            (�(                            ( ��    @           @A       ������������������������������� �(                            (�(                            ( ��    @            @"       �����Ϙ�8�cv?��f?����������� �(                            (�(                            ( �� �q'0g�,���p��s @9<�`  ���u��_��M]u�����u������o��� �(                            (�(                            ( �� �	(�H�(��� %R ��ED�  ���u��_�~�A�����u�����
���� �(                            (�(                            ( �� �y/�H��"�S�xS�� @ED�  ���uv�߷}��_��w����u���������� �(                            (�(                            ( �� ��( H�("�R �	R � @EE  ���uw7_�}�]]��w���u����Ϻ����� �(                            (�(                            ( �� ��ȠH�(��" �%R �@E0E  ����x����c�?��n?�����/�
���� �(                            (�(                            ( �� �x� '�"�!�x��r�8�<�  ����������������������������� �(                            (�(                            ( �� � �                       ������������������������������ �(                            (�(                            ( �� �                    x    ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                      ������������������������o����� �(                            (�(                            ( �� �     �          �    ������������������������o����� �(                            (�(                            ( ��       �          �    ��������?(�ln�lm��~S��)���� �(                            (�(                            ( ��  x�fr��c�����A��p�9�  ������k�}t�kk�k�������w�f����� �(                            (�(                            ( ��  E��� ��@�QTRAA2�"�E   ��������a}�kh?k��������n����� �(                            (�(                            ( ��  E�� ����QTUAA"�"�}   ���������}�kk�k��������n����� �(                            (�(                            ( ��  E"� �� �QTUAA"�"�A   ��������]u�kk������~˾�w�n����� �(                            (�(                            ( ��  E�� ��@dSTH�4A"�"�E   ��������߫l�r�lw(]������� �(                            (�(                            ( ��  x�r T��C����׀�pQ9   ������������������������������� �(                            (�(                            ( ��  @         @              ������������������������������ �(                            (�(                            ( ��  @        �              ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��     P              ������������������������������� �(                            (�(                            ( ��      P  H             ������������������������������� �(                            (�(                            ( ��      P  H             ������?�2�~ڔ�4�6��
�>iƜ��� �(                            (�(                            ( �� �q'0�y�S�%k��y8�c��9c�  ���u��^�u֯�ڳ�}ֺ��k���o���� �(                            (�(                            ( �� �	(� �)PA%L�,�)EE�AY�@  ���u��_u֬>��~|�����.��?��� �(                            (�(                            ( �� �y/���)S�UH���EEA�=�  ���uv�߿u֫���}�}�����뮺���� �(                            (�(                            ( �� ��( @�)TAUH�(�EEAQE@  ���uw7^�u֫�v�}�}ֺ���뮺���� �(                            (�(                            ( �� ��ȡ �)T@�H�(�)EEAQE@  ����x�?�6�?v�~~6��
�>.��/��� �(                            (�(                            ( �� �x� �y�S��(���y8����=�  ����������������������������� �(                            (�(                            ( �� � �           @   @       ���������������������������� �(                            (�(                            ( �� �   �         @  �       ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ���{��������������������������� �(                            (�(                            ( �� �   @           @     ���{��������������������������� �(                            (�(                            ( �� �   @   H              ���{��������������������������� �(                            (�(                            ( �� �   @   H              ���z���ڧ������p��v����� �(                            (�(                            ( �� �d�N%X�k��,��V�    ���zj�[�ښ�]�]mu���뮦������� �(                            (�(                            ( �� ���A%eL����)QYI    ���z���ں�A��mu���.�������� �(                            (�(                            ( �� ��O%EH�"��)��QI    ���z����ں�_��mu������������ �(                            (�(                            ( �� �Q%EH�"��)QI    ���z��[���]�]mu���뮮������� �(                            (�(                            ( �� ��QEH����iQQF    ���������c��m[�p��{����� �(                            (�(                            ( �� y�OD�(����A�Q�    ����������������������������� �(                            (�(                            ( ��            �  �       ����������������������������� �(                            (�(                            ( ��      `�     �          ������������������������������� �(                            (�(                            ( ��                            ������_�����������������￿���� �(                            (�(                            ( ��   �         @    @@   ������������������������������ �(                            (�(                            ( ��   �         @  @  @   ������������������������������ �(                            (�(                            ( ��   �         @  @  @   ����8�T���������j�i������� �(                            (�(                            ( �� y�'�	+','s�@�l�VNX   ���u�WS]��WM�_mu�j�릶������� �(                            (�(                            ( �� �(���	,������AYIYQd   ���t�W]�WW��Xm�������ꮯ����� �(                            (�(                            ( �� ��(��
��"���UAQIQPD   ���u��W]�WW��Wm}�������ꮯ����� �(                            (�(                            ( �� �(��
��"���UAQIQPD   ���u�WW]��W]�Wsu�ھ뮶��n������ �(                            (�(                            ( �� �(���H�����%AQI�QD   ����8�Wa��X���w��ڿn��n������ �(                            (�(                            ( �� y�'��H�"'�r%@�(��ND   ������������������������������� �(                            (�(                            ( ��                         ������������������������������� �(                            (�(                            ( ��     <     0               ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( ��  P    P �            �������������������o���������� �(                            (�(                            ( ��   P $   @�    �       ������������������o���������� �(                            (�(                            ( ��   P $   @� � �       ����2��q��m�N?����&4����
���� �(                            (�(                            ( �� y�S�5�XS���x"��88�`  ���u֯�ٮ��5߀G�]m�}���o��� �(                            (�(                            ( �� �)P@&QdTT� ���,�DE�  ���u֬?۠����t���]m�}������� �(                            (�(                            ( �� �)S�$_DT��`��(�D}  ���u֫�ۯ����u��G�]m�}������� �(                            (�(                            ( �� �)T@$PDT� ���(�DA  ���u֫�ۮ��u߀��Ym�}������� �(                            (�(                            ( �� �)T@$QDTR� x��(�DE  ����6�7뱻�n�v?���7~���
���� �(                            (�(                            ( �� y�S�NDS����Iȁ88�  ������������������������������ �(              �            (�(                            ( ��            �           ����������������������������� �(                            (�(                            ( �� �                     �   ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( �� �                      ������������������������������� �(                            (�(                            ( �� "                    ������������������������������� �(                            (�(                            ( �� "                    ����8�f2T��c*���4�i�g�i������ �(                            (�(                            ( �� "��ͫ��8�c��3�<�`   �����}���]�]j��}�]k���ߦ��o���� �(                            (�(                            ( �� #(�P),����,��Y P YE�   �����~��]�]j����]�.�/�.��o���� �(                            (�(                            ( �� "/��(���<�G��#�E�   ������m��]�]j����]����ۮ��o���� �(                            (�(                            ( �� "( �)(���D�$P$QE�   �����}���]�]j��}�]k���ۮ��o���� �(                            (�(                            ( �� "(�R)(���D�(��QP$QE�   ������vWa�cj���7c�n�7�.�k���� �(                            (�(                            ( �� "'�訞��<Ȝc��#�<�   ������������������������������ �(                            (�(                            ( ��        �                  ������������������������������� �(                            (�(                            ( ��       <                   ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ��                             �/������������������������������/����������������������������� ��                            ������������������������������� �                             �                              ��                            ��                               �?������������������������������?����������������������������� ��                            ��                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ��������������������������������                                ��������������������������������                                ��������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            