�P  �>  P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����                               �����                               �����             �����             �����    �����    �����                       �����    �����             �����    �����    �����                       �����    �����             �����    �����    �����                       �����    �����             �����    �����    �����                       �����    �����             �����       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P - ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    ���       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P ���������                    ���������                              ���������                              ���������                              ���������                              ���������          ������������������          ������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$�I I$�$����O����$�I 	$$�~�������~1$�I#I$�$�1���O����1$�I#	$1$�N�s�ܶ�N�r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1$�I#I$�$�1$�I#	$1$�N s��N r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#O��$�1���I$���1$�I#	$1$�N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#I$�$�1���O����1$�I#	$1$�N s��N r$�I I$�$����O����$�I 	$$�~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$�I I$�$����O����$�I 	$$�~�������~1$�I#I$�$�1���O����1$�I#	$1$�N�s�ܶ�N�r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1$�I#I$�$�1$�I#	$1$�N s��N r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#O��$�1���I$���1$�I#	$1$�N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#I$�$�1���O����1$�I#	$1$�N s��N r$�I I$�$����O����$�I 	$$�~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$��I$�$����O����$�I 	$$�~������~1$��I$�$�1���O����1$�I#	$1$�N�s���N�r���O����$��I$�$�$�I 	$$�~ ��� ~1���O����1$��I$�$�1$�I#	$1$�N s��N r���O����$��I$�$�$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$��O��$���I I$���$��	$$�~ ��� ~1$��O��$�1��I#I$���1$��	$1$�N s��N r$��O��$���I I$���$��	$$�~ ��� ~1$��I$�$�1��I#O����1$��	$1$�N s��N r$��I$�$���I O����$��	$$�~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$�I I$�$����O����$�I 	$$�~�������~1$�I#I$�$�1���O����1$�I#	$1$�N�s�ܶ�N�r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1$�I#I$�$�1$�I#	$1$�N s��N r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#O��$�1���I$���1$�I#	$1$�N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#I$�$�1���O����1$�I#	$1$�N s��N r$�I I$�$����O����$�I 	$$�~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$�I I$������O����$�I 	$$�~������ ~1$�I#I$���1���O����1$�I#	$1$�N�s�ܶ�N r���O����$�I I$���$�I 	$$�~ ��� ~1���O����1$�I#I$���1$�I#	$1$�N s��N r���O����$�I I$���$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$�I O�������I$�$�$�I 	$��~ ��� ~1$�I#O����1���I$�$�1$�I#	$1��N s��N r$�I O�������I$�$�$�I 	$��~ ��� ~1$�I#I$���1���O��$�1$�I#	$1��N s��N r$�I I$������O��$�$�I 	$��~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$�I I$�$����O����$�I 	$$�~�������~1$�I#I$�$�1���O����1$�I#	$1$�N�s�ܶ�N�r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1$�I#I$�$�1$�I#	$1$�N s��N r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#O��$�1���I$���1$�I#	$1$�N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#I$�$�1���O����1$�I#	$1$�N s��N r$�I I$�$����O����$�I 	$$�~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    x  � � x  � �           ���������     @ �       @ �            ��������     @ �  ���O����������~ ��� ~1���O����1���O����1����1��N s��N r$�I I$�$����O����$�I 	$$�~�������~1$�I#I$�$�1���O����1$�I#	$1$�N�s�ܶ�N�r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1$�I#I$�$�1$�I#	$1$�N s��N r���O����$�I I$�$�$�I 	$$�~ ��� ~1���O����1���O����1����1��N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#O��$�1���I$���1$�I#	$1$�N s��N r$�I O��$����I$���$�I 	$$�~ ��� ~1$�I#I$�$�1���O����1$�I#	$1$�N s��N r$�I I$�$����O����$�I 	$$�~ ��� ~���O�������O����������~ ��~ ~x  �$� x  ���      	$   �����������������p  �$�      	$   ����0��p  ��� p  �$�      	$   ��������p �����p �����   ����� ������������UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����