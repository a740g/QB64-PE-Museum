�P  `EO ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                               ��                               ��                               ��                               ��                               ��                               ��                               ��              ����������������@� 0                           �� 0                           �� 0                           �� 0                           @�                             s��                             s��                             s��            ����������������@�                             y��                             y��                             y��                             @�7���                         |��7���                         |��7���                         |��7���        ����������������@����6�                         ~>����6�                         ~>����6�                         ~>����6�                         @�����                         ~>�����                         ~>�����                         ~>�����        ����������������@����3�                         |�����3�                         |�����3�                         |�����3�                         @�0ٶ�6�                         y��0ٶ�6�                         y��0ٶ�6�                         y��0ٶ�6�        ����������������@�0ٶ���                         s��0ٶ���                         s��0ٶ���                         s��0ٶ���                         @�                               ��                               ��                               ��              ����������������@�                               ��                               ��                               ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��  ������������������������     ���  ������������������������     ���  ������������������������     ��                               ����������������������������������������������������������������������������������������������������������                      ����������?���������������������������������?���������������������������������?��������������������������������@                           ����?��������������������������������?��������������������������������?�������������������������������@                           ����?���������������������������������?���������������������������������?��������������������������������@                           ����?���&������g�|8�w��?�������������?���&������g�|8�w��?�������������?���&������g�|8�w��?������������@                           ����?���n��u�ڻۯ���Y��뫿�������������?���n��u�ڻۯ���Y��뫿�������������?���n��u�ڻۯ���Y��뫿������������@                           ����?��]n��u�ڃۯ���[��뫿�������������?��]n��u�ڃۯ���[��뫿�������������?��]n��u�ڃۯ���[��뫿������������@                           ����?��]n��u�ڿۯ�}�[��뫿�������������?��]n��u�ڿۯ�}�[��뫿�������������?��]n��u�ڿۯ�}�[��뫿������������@                           ����?��]o?�u�ڻۯ���[���+�������������?��]o?�u�ڻۯ���[���+�������������?��]o?�u�ڻۯ���[���+������������@                           ����?���o{��W���o�|8k���?�������������?���o{��W���o�|8k���?�������������?���o{��W���o�|8k���?������������@                           ����?����w����������������������������?����w����������������������������?����w���������������������������@                           ����?����������������������������������?����������������������������������?���������������������������������@                           ����?����������������������������������?����������������������������������?���������������������������������@                           ����?����������7����������������������?����������7����������������������?����������7���������������������@                           ����?���}�����������������������������?���}�����������������������������?���}����������������������������@                           ����?���}�����������������������������?���}�����������������������������?���}����������������������������@                           ����?���<8������8�&�1���������������?���<8������8�&�1���������������?���<8������8�&�1��������������@                           ����?��]}�{u�]�5�Z�n�뾦���������������?��]}�{u�]�5�Z�n�뾦���������������?��]}�{u�]�5�Z�n�뾦��������������@                           ����?��]}�{u�]��nn������������������?��]}�{u�]��nn������������������?��]}�{u�]��nn�����������������@                           ����?��]}��u�]���v�n�뮮���������������?��]}��u�]���v�n�뮮���������������?��]}��u�]���v�n�뮮��������������@                           ����?��]}�{u�]���Z�o>뮮���������������?��]}�{u�]���Z�o>뮮���������������?��]}�{u�]���Z�o>뮮��������������@                           ����?��c�8��Wa{�8g�0����������������?��c�8��Wa{�8g�0����������������?��c�8��Wa{�8g�0���������������@                           ����?���������������������������������?���������������������������������?��������������������������������@                           ��  �������������������������������  �������������������������������  ������������������������������   �                           ��  ������������������������     ���  ������������������������     ���  ������������������������     ����                       ����������������������������������     �����������������������������     �����������������������������     ��                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          ������������������������������������������  ������������������������������������������������������������������                      ������������������������������������������������������������������                      w�����{���������������w�����{���������������w�����{���������������                      �����{��������������������{��������������������{���������������                      ~2m��+N18����L�c���`~2m��+N18����L�c���`~2m��+N18����L�c���`                      ������j�7��}���5��w�頍�����j�7��}���5��w�頍�����j�7��}���5��w��                      �����jv�}���u��w�������jv�}���u��w�������jv�}���u��w��                      ������j�u������u��w��������j�u������u��w��������j�u������u��w��                      u�����j�u��~n��u��w��u�����j�u��~n��u��w��u�����j�u��~n��u��w��                      �6���kv�����v�ㇳ렎6���kv�����v�ㇳ렎6���kv�����v�ㇳ�                      ���������������������������������������������������������������                      ������������������������������������������������������������������                      ������������������������������������������������������������������                      �����������o�������������������o�������������������o��������                      ���������������������������������������������������������������                      ���������������������������������������������������������������                      vq���N3����q�>M�8cS�vq���N3����q�>M�8cS�vq���N3����q�>M�8cS�                      u��m���5�ڻ�k���ݿ�}M�u��m���5�ڻ�k���ݿ�}M�u��m���5�ڻ�k���ݿ�}M�                      v��m��tڃ��0�ݾa]�v��m��tڃ��0�ݾa]�v��m��tڃ��0�ݾa]�                      wo�m��u�ڿ�����ݽ�]]�wo�m��u�ڿ�����ݽ�]]�wo�m��u�ڿ�����ݽ�]]�                      e��s��u�ڻ�뮵��}�]]�e��s��u�ڻ�뮵��}�]]�e��s��u�ڻ�뮵��}�]]�                      �q���v7����p�?^�a]`�q���v7����p�?^�a]`�q���v7����p�?^�a]`                      ���������������������������������������������������������������                      ������������������������������������������������������������������                      ������������������������������������������������������������������                                                �  ������������������������������������������������������������������                      �?���������������{�����?���������������{�����?���������������{����                      ���������������������������������������������������������������                      ���������������������������������������������������������������                      ��ɷ�|�~���8]�f8{>�g���ɷ�|�~���8]�f8{>�g���ɷ�|�~���8]�f8{>�g�                      �7[��k����]��]u��z�k���7[��k����]��]u��z�k���7[��k����]��]u��z�k��                      ��[���=�>�]�]�{~����[���=�>�]�]�{~����[���=�>�]�]�{~��                      ��[�������]��]m�{�����[�������]��]m�{�����[�������]��]m�{���                      ��[��뽫�7Y��Yu��z�����[��뽫�7Y��Yu��z�����[��뽫�7Y��Yu��z���                      �8����}�x��8e�v8{>�w��8����}�x��8e�v8{>�w��8����}�x��8e�v8{>�w�                      ������������������������������������������������������������                      ���?��������������������?��������������������?�����������������                      ������������������������������������������������������������������                      ������������������W���������������������W���������������������W���                      ���������������������������������������������������������������                      �����������߯�������������������߯�������������������߯��������                      �>�8�o1�8Ɏ��'^V?���>�8�o1�8Ɏ��'^V?���>�8�o1�8Ɏ��'^V?��                      ���u�[on��[u�vj��^�������u�[on��[u�vj��^�������u�[on��[u�vj��^����                      ��u�[on��[�v��������u�[on��[�v��������u�[on��[�v������                      ���u��on��[}������������u��on��[}������������u��on��[}���������                      ���u�[�n��[u�����~�������u�[�n��[u�����~�������u�[�n��[u�����~����                      ��8ۿq��m����^�7����8ۿq��m����^�7����8ۿq��m����^�7��                      ������������������������������������������������������������������                      ���������������������������������������������������������������                      ������������������������������������������������������������������                      ������                    �  ������������������������������������������������������������������                      ���������������������������������������������������������                      z�������������������z�������������������z�������������������                      z�������������������z�������������������z�������������������                      z�����N?�ƙm�q�<�`z�����N?�ƙm�q�<�`z�����N?�ƙm�q�<�`                      ��]���{5�뭺km뾺뽫���]���{5�뭺km뾺뽫���]���{5�뭺km뾺뽫�                      ~�����{t����m밺�� ~�����{t����m밺�� ~�����{t����m밺��                       ~����v��u�����m뮺����~����v��u�����m뮺����~����v��u�����m뮺����                      ~��]�ww{u��-��s뮺뽫�~��]�ww{u��-��s뮺뽫�~��]�ww{u��-��s뮺뽫�                      ~���x�v?���w�p�=�`~���x�v?���w�p�=�`~���x�v?���w�p�=�`                      ������������������������������������������������������������������                      ������������������������������������������������������������������                      ������������������������������������������������������������������                      ���������������������������������������������������������������                      ���������������������������������������������������������������                      ���������������������������������������������������������������                      �������~f3c�8|1����������~f3c�8|1����������~f3c�8|1���                      u������[~���]���{����u������[~���]���{����u������[~���]���{����                      u�����PU~�-�]���{����u�����PU~�-�]���{����u�����PU~�-�]���{����                      u�������~����]u��{����u�������~����]u��{����u�������~����]u��{����                      u������n����]u��{����u������n����]u��{����u������n����]u��{����                      ��������n7c��|1�����������n7c��|1�����������n7c��|1���                      ���������������������������������������������������������������                      ������������������������������������������������������������������                      ������������������������������������������������������������������                      ����������������          