�P   ˀ�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ������������������������������������������������������������������������������                                                                                                                                                                                                                                                 �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �������������������������������������������������������                        ������������������������������������������������������                                                                                                                                                                                        ������}��������}�����ٻ���������������������������                           �   P@ ��  �@ H�   (P  � � ��   �                                                                                                            @�     �  &D "  �B  �   $ �@@ (�D                        �������������^�����}�����v�������������_o������������(                         @��  ��@!�@` �      � � B   (	  � 
                                                                                                           	    �	   � $ (�  @�@B 	  ��         �                        �}���������߯}��߿��}�6����}���w���������������������                        1 @ �     D$de    �    PH A   D �                                                                                                           �   @  P�  @��� �p " �  �@D @  	 A   $                        ����������o�v�����������������y��������������a�����                          �     @A A �X��  ��!(  !@�  @�   �                                                                                                             � �S D� �   �          �@ h@ @ � �QB                        ��?���������{~���������������?�W���������a�=�����������                          @   � @  "  � �   @ P�        �    ��                                                                                                          D�  @P	�� @%   ! "  �0�     � �hP@   P  L                        ��_�������~����������������_����ޗU���������|��������0                        �  @��       @ @1PPH T       @ �  @@                                                                                                          *�   �     `  �  0	!h�   d$H �  !  �                        ������������������������������������������o�����~��                        <�(  D d@ 
 K� H0   �P ���I   D	!@$ A  Ԅ BH                                                                                                          B0  (�   �   �!      �0   �  �                        ��}����������������_�?��������=����7�������g�������                         P1  �E@ h@ !      A  � � ` (@ �                                                                                                           A�  �       �� �B!  DC  �(�   @ �                             ��_߿���������������������_�?�������g�������������}}�                          �B $	       B� 
 �  \�H �  *  H @                                                                                                             � @    H�! D     @� �     �         ��                        ���                                                  �                        �                                                   `                                                                                                           ���������������������������������������������������                        �����������������������������������������������������x                         ?���������������������������������������������������                            ?���������������������������������������������������                           @                                                  �                        �ݿ����������������������������������������������������                        ?���������������������������������������������������                            ?���������������������������������������������������                           "@                                                  $                        ���                                                  ��                         ?���������������������������������������������������                            ?���������������������������������������������������                            O��������������������������������������������������                         ��7����������������������������������������������������                        �8                                                  �P                           ?���������������������������������������������������                            ���������������������������������������������������                         ��7����������������������������������������������������                        �8           @                     @          ��                           ?���������������������������������������������������                            ���������������������������������������������������                         ��7������������������������������������������                        #8 ���}����cA��������4 ���}����cA��������4�0                           ?�������     �������     �������     �������     �                           @�     �     �     8          �     �     8                             ������>���w�|��������������>���w�|�������������                         8  ��������@ �������84  x��������@ �������84�                            ?�������     �������     �������     �������     �                           N     �     �     8         �     �     8      t                        ������ ����e����������[����� ����e����������[���x                        `8 ��}����#@��������4 x��}����#@��������4�                            ?�������     �������     �������     �������     �                           N     �     �     8         �     �     8      �                        ������������\�����8��������?�����\�����8������x                        @9���������X��������5��?������X��������4�                            ?�������     �������     ���?���     �������     �                           N     �     �     8       ?� �     �     8      �                        ��������ꏾ������>���8|�[��� �ꏾ������>���8|�Z��                         9�������x4�\������O���?����x4�\������O��                            ?�������     �������     ���?���     �������     �                           N     �     �     8       ?� �     �     8      d                        ��������������?(�����;������������?(�����:��                         9������x4�\8��������O�������x4�\8��������O��                            ?�������     �������     �������     �������     �                           �N     �     �     8         �     �     8                             �߶��~��~���_H�����-����q���x��~���_H�����-����u���                        9����?�߸��\ 9������}�����?�߸��\ 9�������}��                           ?�������     �������    �������     �������     �                            N     �     �     8        �     �     8                             �ζ/���o������������O��A�/��o������������O���A���                         9��������_�`_�п����5��������_�`_�п����4�                            ?�������     �������     ������     �������     �                           1N     �     �     8  >    � �     �     8                             �������������P��������`E���������P����������E
��                        P9� ��A����_� ����`������A����_� ���������                            ?�������     ������� 0 ������     �������     �                            N     �     �     8 ��  �� �     �     8                              ����������S�?�����(�� C���  ���S?�?�����(��7�C���                        ������q�����_�+@��� ��   ��q��?��_�+ �������                           ?�������     ������� D ��  ���  �  �������     �                            N     �     �  p  8 ��  �� � �  �     8                              ����������~������h��  G���  ���~������h��y�G���                        �9�����s����_�~��?� ���  ��s��?��_�~8��?�����                            ?�������     �������     ��  ���     �������     �                           N     �     �  p  8 ��  �� � �  �     8                             �����?���O��?���/��  z� ?�����?����/���� z��                         9���� �����_���� ���  �� ����_�<��������                            ?�������     �������     �� ���    �������     �                           �N     �     �  �  8 ��  �� � �  �     8                             ���}�q����?_����c���� �| ����9��������������X                         9�����_����_�p`�Pu� ���� ��_����_�p(�Pu������                            ?������     ���S���     �� ��� @  ������� >8 �                           ZN �� �     � �  8 ��  �� � �  �     8 >8 �                        ��=�pw���@����A��  !�> w���A�������&�!���                         ����������_l@�Pp� 	���� �����_c��Pp������                           ?��p}���     ���9���     �� ���  �  �������  0 �                           �N �� � 0   � �  8 ��  �� � �  �    8 >8                         �z�̽�p'��� ?�>������  c�̿ '���8�>���?�����c���                        h9����s/����_�� �W2� ���� �s/���_��0�W2������                           ?��p}���     ���1���     �� ���  �  ���?���  0 �                           �N �� �    � �  8 ��   �� � �  � �  8 >8 T                        ������ o��C��>�� ����< C��� o��C��>�����7�C���                         9����w� ��[����W{� ���� �w���[���W{�����                            ?�� }���    �������     �� ���    ������ � �                            N �� � �  �   8 ��   �� � �  � �  8 ��                          �?�������A�f�� @����� Fk�  ������f��A�����  Fj��                        "9����e�A��\_�@�W�  ���� �e���\_�@�W� ���                            ?��0��� �  �������     �� ���    ������� �p �                           �N �� � ��  � �  8 ��  �� � �  � ?�  8 ��                         ���������  y��� ���������������d y��� ���� ����                         8	� �� ��@� ������t� �����@� a��� �t�                            ?��0��� @   �������   �������    ����� �p �                           N �� � ��  � �  8 ��  �� � |  � ?�� 8 �� $                        ��������  ��������� ����  ���� ���� ?���� ����                         8� ��  �@ ���� �4   ���C�@   ��� �4�                            ?��0��� �  �������     ��  ��� �  ���?�� �p �                           �N �� ���  � �  8 ��  �� � �  � �� 8 ��                         ���������  ~>��� ��o�������� ��� ~>��� ?�o�� ����                        	8� ��  ��@  ������� �����@   ��� ��                           ?��0��� 0   ������ > ����  @  ��� ?�� �p �                            N �� ���  � �  8 ?��  ���� �  � �� 8 ��                          ���������� ���� ?�)�� ����  �������  �)�� ����                        �9�� ��� �X ���� ��   ��� ��X   ��� ��                            ?��0��� `  ������     ��  ���     �� ��� �p �                           `N �� ���� � �  8 ��  �� � �  � ��� 8 ��                         ��������� ?����?��� 7�����������0 ��� ����                        ����  ��� ?�_� ��?� O�e�   �����_�0  �?� �d�                           ?��0���     ������     ������     ��  �� �p �                           N �� ���� � �  8  ��   ?� � �  � ��� 8 ��  $                        ���� �ҽ�  ?�����+�� �����ҽ�� ��@ �+�� ����                        ��   }C�  ?�_� ��?� �E�   }C����_�@  �?� �D��                           ?�� ���   ������     ������     �� �O��     �                            N �� ���� � �  8  ��   ?� � �  ���� 8 ��                          ���������  ?������� �K������� ��� ��� �J��                         9�   mG�  ?�_� ��� ���   mG����_��  �� ?���                            ?������   ������     ������     �� �O��     �                            N  � ���� �  �  8  ��   ?� � �  ���� 8 ��                          ����������  �������� ��������� ���  ��� ����                         9�   g�  �_  � V� ���   g����_    V� ���                            ?������    ������     ������     �� ���     �                           @N  ?� ���� � �  8  ��   ?� � �  ���� 8  ��                         ��7�� ����  �����?��� ���������� ���  ��� ����                        8�   �  �N �  �� ?���   �� ��N     �� ���@                           ?�� ��� � � ���8?��     ������ �  ��  '��     �                            � �� ���� � �� 8 ��   � � �  ���� 8 ��                         ����� ����  ���� ���� ���������  ���  ���� ����                        �8     �  �@     �� ?��    �  �@     �� ����                           ?�� ��� B � ��� ��     ������     ���'��     �                            N �� ���� � ?�� 8 ��   � � ��� ���� 8 ��                          ������ ����  ��� ���� 6��������< !��  �������                        E8 � ~�  �@  ��� ?��   ~�< >�@  ������P                           ?������ � ������     ������ 3�� ��- '�� x �                            N �� ���� � �� 8 ��   � ���� ���� 8 ��                          ���� ����  ?��� ���� 6��������  a?�� ���� ���                        (8    �  �@   ��� ?��   �  ~�@   ��� ���                           ?�� ����   ��� ��     ������     ��: ��     �                           N �� ���� � ?�� 8 ��   � � ��� ���� 8 ��                         �Ƿ���?����@  ?�������� ��� ������?�� ��������x                        B8    �@ ?�@   ��� ��    ����@   ��������                            ?���?����   ������     �� ���     ��4 ��     �                           8N  � ���� � �  8 ��   �� � �  ���� 8    �                        ������?����� 0�������� ��� �����p��  ���������                        �8   ?��� ?�@   #��� ��   ?�����@   ��������@                           ?���?���   ������     �� ���     ��h O��     �                           AN  � ��� � �  8 ��   �� � �  ���� 8                            ������?����@ �������� ���� ����� ���� ���������                         �   <��@ �@  �8�� ��   �����@   8�������                           ?���?���    ������     �� ���     ��� ���     �                           N  � � ��� � �  8 ��   �� � �  � ?�� 8     d                        ���������� ?��������� ���� ��������� ���� g����                        8@   �� ?�D   ` �� ��@   ����D     �� ���                           ?������ @   ������     �� ���     ��� ��     �                           �N  ?� ���� � �  8 ��   �� � �  � �� 8  ��                         ����������@ ��������������x���������� ���� {����                        �    �@ �@    �����  x ����@    �� ����                           ?������ � @ ������   ��G���     ��� ��     �                           N  ?� ���� � �  8 ��  �� � �  � �� 8  ��  t                        ��������?  ?���� ��������������?������ ���� ;����                         8   �  ?�@p   ����� � ����@p    �� ?���                            ?������  � ��� ��� � ������     ��� o��     �                           �N  � � ��� � �  8 ��  �� � �  � ?�� 8 ��                         �۷�������~ ?���� ���������� �������������� ;����                         ���  ~>~ ?�[�   ���������  ~?���[��  ��� ?���                           ?������ a�  ��� ���   ������     ���|��     �                           $N  � ���� � �  8 ��  �� � �  � �� 8 �� D                        ���������  ���� ��������� ���������� ��� 9����                        "9�� �~?  �]�   ������� �~?���]�   �� ?���                            ?������     ��� ��� 
@ ������     ��� ��     �                           N  � � ��� � �  8 ��  �� � �  � ?�� 8 ��                         ��7�<����� ��������� ���x� ����� ��������������                        9��< ���X��P �� �����  ���X��P ������@                           ?��#���� 	�  ���p�� � �� ��� 	�  ���p��  �  �                            �  �� � ?�  � �� 8 ��  �� � ?�  � �� 8 ��                         ��7��p���?� ���� ?���� ����  ���?� ���� ?���������                        8 p �� ��@p   �� ��    �� ��@p   ������                           ?��H���   ��� ���    �� ���   ��怿��    �                           @� �� � �  � �� 8 ��  �� � �  � �� 8 ��                         ���������< ���� ���� ����  ��� ���� ���������                        � �  �< �@    W�� ��    �� �@    W�������                           ?������ 2  ���_��    ��  ��� >  ��̀_�� � �                            N �� � ��� � �� 8 ?��  ���� �� � ?�� 8 ��                          ����������8 x���� ���  ���  ���< x���� ���3��
��                        �8�� �8 �@ ���� ���  �< �@ ��������                            ?��L���  � ��Ā?��     ��  ���  � ����?�� 0 �                           `N �� � ��� � ?�� 8 ?��  ���� ��� � ?�� 8 ��                         �߷� ����  y��� ���  ���   ?���  y��� ��� ����                        A8�  x  �G�� �׀   ���  x  �G�� �׀p ���                           ?������ < � ��� ?��    ��  �� < � ��� ?�� � �                            N �� � ��� � ?�� 8 ��  ���� ��� � ?�� 8 ��                         �߷    ����  ?��   ���� � � ���  ?��   ���� ����                        �9��   @   ?�_��   � � ����  @   ?�_��   �   ���                            ?�� ���   @ ��� �� x�����?��   @ ��� ��    �                            N �� ���� � �� 8 ���� ?������� � �� 8 ��                         ���    ����  ?��   ���   �    ���  ?��   ���� ����                        9��       ?�_��       ���       ?�_��      ���                            ?�� ���   @ ��� ��    ���  ?��   @ ��� ��    �                            N �� ���� � �� 8 ���� ?������� � �� 8 ��                          ����� ?���� �� � ���   ��   ���� �� � ����� ����                        9���   � �_��       ���    � �_��    � ���@                           ?�� ���� ������    ���  ?���� ������ | �                            N ������� ���� 8 ���� ?������� ���� 8 ��                          ��7�   ?���  ��   ���   ��   ���  ��   ����  ����                        9�   p   �W�        ��   p   �W�        ���                            ?��  ��    ��  ��    ���  ?��    ��  ��    �                            � ������� ���� 8 ���� ?������� ���� 8 ��                          �߶�   ?���  ���  ��   ��   ���  ���  �쟀  ����                         9��   6   �_�    `   ���   6   �_�    `   ���                            ?��  ��    ��  ��    ���  ?��    ��  ��    �                            N ������� ���� 8 ���� ?������� ���� 8 ��                         �������������������������������������������������������                         8           @                     @          �                            ?���������������������������������������������������                            O��������������������������������������������������                         �ִ                                                 �h                         ;���������������������������������������������������                            ?���������������������������������������������������                           )O���������������������������������������������������                        �������������������������������������������������������                        �8           @                     @          �                            ?���������������������������������������������������                            O��������������������������������������������������                         ������������c��!��/����;���������c��!��/����:��                         9����� ?x�_�����`��������� ?x�_�����`�����                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                              ������������������]�/����8;���������������]�/����8:��                        9���>  ��_������ �������>  ��_������ ������                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��������������#���Yo�/����;�����������#���Yo�/����:��                        ���� � @��_������������ � @��_�����������                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      T                        �]�~� }r������`�/����:~� }r������`�/����:��                        �������`A����_����8�����������`A����_����8�������                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     
$                        �=�>�,���x4������o���O�>�,���x4������o���O���                        9������pA����_���>�����������pA����_���>������@                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     $                        ���>�r�,N���x4����/�������O�>�r�,N���x4����/�������O���                        �9������p@����_���?<��������p@����_���?<���                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ���?��}#��߸�߳����>+����}�?��}#��߸�߳����>+����}��x                        8��~��}p x��'O���-�� ��t��~��}p x��'O���-�� ��t�0                           >     �������     ?������     �������     ?�������                           XN     �     �     8          �     �     8     �                        �������r������?��(�����;����r������?��(�����:��                        �/���o��E�B�������W��/���o��E�B�������W���                           >     �������     ?������     �������     ?�������                           cN     �     �     8          �     �     8     4                        �U�����QB����믯���,���������QB����믯���,������X                         9�����  �P������  �������  �P������  ���                            >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     
�                        �;6;�M�P�����������������
;�M�P�����������������
�                         9����� ���\�����
�������� ���\�����
����                            >     �������     ?������     �������     ?�������                           ��     �     �     8          �     �     8     L                        ���38x�������3���?����38x�������3���?������                        9�����1����\�����W���������1����\�����W�����@                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              �����>���������������������>��������������������                         8���?��@��@?����������?��@��@?��������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8     D                        �׷���~ z�_�����/����u��������~ z�_�����/����u������x                        8��������A�������
���������A�������
��@                           >     �������     ?������     �������     ?�������                           (N     �     �     8          �     �     8     �                        �������z�����������p���������z�����������p�������                         8?��w�}����A���������?��w�}����A����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        ��3@�����/�����4���2�?���3@�����/�����4���2�?�����                         9̿�'�����\���������̿�'�����\����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                             ��6a�����������{�?���a�����������{�?�����                         9���o�o����]� �����������o�o����]� ���������                            >     �������     ?������     �������     ?�������                           �     �     �     8          �     �     8      l                        ���;��~������������ >��;��~������������ >���x                         9� ���q���_� ���������� ���q���_� ����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      �                        ������q�n�������XF����?�{���q�n�������XF����?�z��                         9������ B����_������)��������� B����_������)����                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      T                        �����q������������o���?�;���q������������o���?�:�x                        $9����� @��_�������������� @��_����������@                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8     �                        �����1�����������������?����1�����������������?���                        �9����� @ ?��_�����P ������� @ ?��_�����P ����                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                             �;�~�������8�������������
~�������8�������������
�                        9�����`@ ?�_���?� �������`@ ?�_���?� ����                           >    �������  `  ?������    �������  `  ?�������                           �N    � �  �  p  8        � �  �  p  8    D                        �߷��������ƿ� ��h?����k��������ƿ� ��h?����j��                        �8��s�~  �?@��?�� ����s�~  �?@��?�� ���                            >    ������  �  ?������    ������  �  ?�������                            N  � � �  �  �  8  >    � � �  �  �  8  >                          �������������������?����J����������������?����J��                        �9��?��~ ��P������ 8����?��~ ��P������ 8���                            >    ������ �  ?������    ������ �  ?�������                           N  � � �  � �  8      � � �  � �  8     D                        �����������������,�8����������������,�8����                        9����~ ��Q������� 8x�����~ ��Q������� 8x��                            >  -  ���G��� �  ?�����  -  ���G��� �  ?������                            N  ?� � �  � �  8  ��   ?� � �  � �  8  ��                          ���o����������������0��o����������������0����                        9�����| �Y������� 0x �����| �Y������� 0x �@                           >  #  ������� 2  ?������  #  ������� 2  ?�������                            N  ?� � �  � �  8  ��   ?� � �  � �  8  ��                          �w������������� ���� �������������� ���� ���x                        2������8  � _����Ӏ  x �����8  � _����Ӏ  x �(                           >  .  ������� �  ?������  .  ������� �  ?�������                           �N  ?� � �  � �  8  ��   ?� � �  � �  8  �� �                        �77������������� ��������������������� ���������p                         9���?��   � _�����   � ���?��   � _�����   � �                            >  @ ������   ?������  @ ������   ?�������                           ��  � � �  � �  8      � � �  � �  8    �                        �����=�����������_����������=�����������_��������x                        9���?��    ��_�����   	����?��    ��_�����   	��                           >  � ���?���   ?������  � ���?���   ?�������                           N  � � �  � �  8      � � �  � �  8    �                        �w����������?�������O����������������?�������O��������x                        �������    ��_������   	�������    ��_������   	��x                           >    ���?���  @  ?������    ���?���  @  ?�������                           �N    � �  �  p  8        � �  �  p  8    �                        ���������������� ���� ?��������������� ���� ?����                        9�����    �_�� ���   ������    �_�� ���   ���                           >     ������     ?�� ?��     ������     ?�� ?���                           N  � � �  � �  8 ��   � � �  � �  8 ��  D                        �����|�~���������\��������|�~���������\��������                        9��|��   ��_����� ����|��   ��_����� ����                           >  c� ������� <  ?�����  c� ������� <  ?������                           AN  �� � ?�  � �� 8 ��   �� � ?�  � �� 8 ��                         ��7����~�������� ?���� ?������~�������� ?���� ?����                        @9�����    �_�� ���   0�����    �_�� ���   0�                            >     ������     ?�� ?��     ������     ?�� ?���                           �  � � �  � �  8 ��   � � �  � �  8 ��  L                        ������������?������������������������?�����������������                        9������  � _������  � ������  � _������  � ��                           >     ���?���     ?������     ���?���     ?�������                           N    � �  �  p  8        � �  �  p  8     D                        ��7���>����������������������>���������������������                        �9�����   @ _�����   �����   @ _�����   �                            >     ������     ?������     ������     ?�������                            �  � � �  �  �  8  >    � � �  �  �  8  >                           ������~����������������������~��������������������H                        �������  @ _�����   ������  @ _�����   �H                           >     ������     ?������     ������     ?�������                           N  � � �  �  �  8  >    � � �  �  �  8  >   �                        ���G?�>���?����s���/������G?�>���?����s���/��������                        @9���?��o�  @_������   5���?��o�  @_������   4�                            >     ������     ?������     ������     ?�������                           N  � � �  � �  8      � � �  � �  8     D                        ���'?���?����s������ ��'?���?����s������ ����                        49�����w�  ` _�����   �����w�  ` _�����   �@                           >     ������     ?�� ��     ������     ?�� ���                            N  ?� � �  � �  8  ��   ?� � �  � �  8  ��                          ��6s��
�������;�������p?��s��
�������;�������p?����                        9����c�@ _������? p ����c�@ _������? p �@                           >  � ������� 8  ?��N?��  � ������� 8  ?��N?���                           �  � � �  � �  8 ��   � � �  � �  8 ��                         �}���0���������� _���������0���������� _���������                         9��0��� � _�� �� � ��0��� � _�� �� � �                            >  ( ������ �  ?���_��  ( ������ �  ?���_���                           �N  �� � ?�  � �� 8 ��   �� � ?�  � �� 8 �� $                        ��7��p����� ����� ?���������p����� ����� ?���������                        9��p�� �  _�� ?���  ��p�� �  _�� ?���  �@                           >  | ������ �� ?���/��  | ������ �� ?���/���                           � �� � �  � �� 8 ��  �� � �  � �� 8 ��                         ����p��� ����� > /������p��� ����� > /�������                         9��p��� _�� ?���� w���p��� _�� ?���� w��                            >  , ������ �@ ?�����  , ������ �@ ?������                            N �� � �  � �� 8 ��  �� � �  � �� 8 ��                          ���� ���� ����  >~/�x ���� ���� ����  >~/�x ����                         �� ���� ^� ?����  `u� ���� ^� ?����  `t�                           >  x ������ �@ ?�����  x ������ �@ ?������                           �N �� � �  � �� 8 ��  �� � �  � �� 8 ��                         ����� ���   ���� �,   ���� ���   ���� �,   ����                        (9   ���   P   ����   5   ���   P   ����   4�                           >    ��  ���     ?�� ��    ��  ���     ?�� ���                           N �� � ��� � ?�� 8 ��  �� � ��� � ?�� 8 ��  D                        ����� ���   ���� ��   ���� ���   ���� ��   ����                         8   ���    @   ����      ���    @   ����   �                            >    ��  ���     ?�� ��    ��  ���     ?�� ���                            N �� � ��� � ?�� 8 ��  �� � ��� � ?�� 8 ��                          �߷�� ��� ���~ �� ����� ��� ���~ �� �����                         ��� ���   H ~ ���߀  �� ���   H ~ ���߀  �                           >  �����?�� q� ?��|��  �����?�� q� ?��|���                            N ������� � ��� 8 ?��  ������� � ��� 8 ?��                         �����  ��   ���  ��   ����  ��   ���  ��   ����                        9�   �_�    \   ����   �   �_�    \   ����   �                           >    ���  ?��    ?�� ��    ���  ?��    ?�� ���                           @N ������� � ��� 8 ?��  ������� � ��� 8 ?��                         ���'�  ��   ��  ��`  ��'�  ��   ��  ��`  ����                        d��   ��    M�  ����   �   ��    M�  ����   �H                           >    ���  ?��    ?�� ��    ���  ?��    ?�� ���                            N ������� � ��� 8 ?��  ������� � ��� 8 ?��                          �����������������������������������������������������8                         8           @                     @          �                            ?���������������������������������������������������                           O�������������������������������������������������� �                        ���                                                 ��                         ;���������������������������������������������������                            ?���������������������������������������������������                           O�������������������������������������������������� D                        �������������������������������������������������������                        ��           @                     @          ��                           ?���������������������������������������������������                           @O��������������������������������������������������                        ���������������������������������������������                        � ���}����cA��������4 ���}����cA��������4�                           ?�������     �������     �������     �������     �                           pN     �     �     8          �     �     8                             �۷���>���w�|��������������>���w�|�������������                        8  ��������@ �������84  ��������@ �������84��                           ?�������     �������     �������     �������     �                           $N     �     �     8          �     �     8     D                        �Ϸ��� ����e����������[����� ����e����������[����                        8 ��}����#@��������4 ��}����#@��������4�0                           ?�������     �������     �������     �������     �                           0N     �     �     8          �     �     8                             ������������\�����8��������������\�����8������x                        @9���������X��������5���������X��������4�                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        �޷�����ꏾ������>���8|�[�����ꏾ������>���8|�Z��                        �9�������x4�\������O��������x4�\������O��                            ?�������     �������     �������     �������     �                           !N     �     �     8          �     �     8                             ���������������?(�����;������������?(�����:��                        �9������x4�\8��������O�������x4�\8��������O��                           ?�������     �������     �������     �������     �                           dN     �     �     8          �     �     8     D                        �����~��~���_H�����-����u���~��~���_H�����-����u���                        @9����?�߸��\ 9�������}�����?�߸��\ 9�������}��                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ���/���o������������O���A�/���o������������O���A���                        �9��������_�`_�п����5��������_�`_�п����4�                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �������������P����������E����������P����������E
��                        C9� ��A����_� ��������� ��A����_� ���������0                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ����������S�?�����(��7�C��������S�?�����(��7�C���                        9����q�����_�+ ����������q�����_�+ �������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �����������~������h��y�G���������~������h��y�G���                         9�����s����_�~8��?���������s����_�~8��?�����                            ?�������     �������     �������     �������     �                           PN     �     �     8          �     �     8                             �o����?���O��?����/���� z���?���O��?����/���� z��                         9���� �����_�<����������� �����_�<��������                            ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8     	                        �}�������?_������������������?_��������������                         9�����_����_�p(�Pu����������_����_�p(�Pu������                            ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8     $                        ���?��w���@�������$�!�?��w���@�������$�!���                        �9���������_o��Pp��������������_o��Pp������@                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ���̿�'���<?�>���������c�̿�'���<?�>���������c��x                         9����s/����_����W2�?�������s/����_����W2�?����                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        ������o��C�o�>�� ����?��C����o��C�o�>�� ����?��C��x                        9���A�w����[����W{�?������A�w����[����W{�?����                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        ���� ������_�f�� ��������Fk� ������_�f�� ��������Fj��                        �9�����e����\_���W� >�������e����\_���W� >���                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      D                        �߷��������`y���������Ǒ���������`y���������Ǒ���                         8
�������@�������?�t
�������@�������?�t�                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                             ��7������������������9���������������������9�����                        J8 q������@�����?�4 q������@�����?�4��                           ?�������     �������     �������     �������     �                           $�     �     �     8          �     �     8     L                        ������������~>������o���������������~>������o��������                        h8  �������@ �����?�  �������@ �����?���                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �����������������?�)���w����������������?�)���w����                         9�  �������X ��������  �������X ��������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��6�������������?����7���������������?����7���p                        9�  ~ ������_� ��?����e�  ~ ������_� ��?����d�@                           ?�������     �������     �������     �������     �                           �     �     �     8          �     �     8      �                        ������ҽ���������+���������ҽ���������+�������                         9�  ~ }C�����_� ��?����E�  ~ }C�����_� ��?����D�                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                             ���������������������K�������������������J��                        (9�  � mG�����_� ��������  � mG�����_� ��������                           ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8                             ��7���������������������������������������������                        	9�  � g�����_  � V������  � g�����_  � V������                           ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                             ������������������������������������������������x                         8�  ~ �����N  � �������  ~ �����N  � �������                            ?�������     �������     �������     �������     �                           XN     �     �     8          �     �     8     �                        ���������������������������������������������������                        	8   ~ �����@  � ������   ~ �����@  � �������                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �������������a����������������������a��������������                         8  ~�����@  '�������  ~�����@  '��������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �������������a?����������������������a?��������������                        8   �����@   '�������   �����@   '��������@                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    