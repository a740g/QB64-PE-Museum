�P  �>  P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��       ��       ��                 �        �        �                                                                                                                                                                                                                         By��                                 B�D                                 B�D                       �{���    �����                        @ DH    ~�G�H                       @ DH    F�DTH                       �{���    �����                       @ DH    F�DTH                         H    F|G�H             >     |  >�����|  >�����|                     >DDDDH|  >DDDDH|                      >DDDD@|  >DDDDH|                 8   >�����|  >�����|                     >�����|  >�����|                     >�����|  >�����|                     >�����|  >�����|                     >�����|  >�����|                                 �����        �����                     ]����       �����       �����                     �����       �����       �����                    �����       �����       �P - ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������� �������� �������� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������/��������/��������/��������/�������{���������{���������{���������{���������{���������{���������{���������{��������    7�����    7�����    7�����    7������;�+�������;�+�������;�+�������;�+�������;���������;���������;���������;��������    7�����    7�����    7�����    7������;���������;���������;���������;����������� ��������� ��������� ��������� ������    7�����    7�����    7�����    7�������������������������������������������������������������������������������������    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    ���~��?���  ?����������  ?�~��?���               >0f��3`��  ?����������  ?�~��?���               ?�~��?���  ?����������  ?�~��?���               >0f��3`��  ?����������  ?�~��?���    P                               ������������������������������������          ���������������������������          ���������������������������                    ������������������          s��9�s��9�������������������          ���������s��9�s��9�s��9�s��9�          c�1�c�0���������s��9�s��9�          ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              o���������������� ����           }k�����_־�8p�9��8p�9�          o�������~��/�_���~�(
P�)@          ���������b��#F b��#F           ���������������������?��          ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           |����>���?�� @           |����>��������� @           |����>���?�� @           ���������������������?��          ��������� @  @           |����>��������� @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           |����>���?�� @           p ��� p ���           ��?���������������?������?����          p ��� �����������?����          ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           |�����>��������� @           |�����>��?��� @           |�����>��������� @           ������������?�����?��          ���������|����> @           |�����>��?��� @           |�����>��������� @           |�����>��?��� @           |�����>��������� @           |�����>��?��� @           |�����>��������� @           p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                                                  ������������������������������������          ���������������������������          ���������������������������                    ������������������          s��9�s��9�������������������          ���������s��9�s��9�s��9�s��9�          c�1�c�0���������s��9�s��9�          ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           |����>��������� @           |����>���?�� @           |����>��������� @           ������������?�����?��          ���������|����> @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           �������|������> �          ��������?�@  �          �������|������> �          ����������?���?��          ���������|����> @           ��������?�@  �          �������|������> �          ����������?�@ �� �          |�������������> ���      |��������?�@  �          |�������������> �          p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           |����>��������� @           |����>���?�� @           |����>��������� @           ������������?�����?��          ���������|����> @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           |������>��������?�@           |������>�� ��?�@           |������>��������?�@           ������������?�����?��          ���������|����> @           |������>�� ��?�@           |������>��������?�@           |������>�� ��?�@           |������>��������?�@           |������>�� ��?�@           |������>��������?�@           p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           |�����>�������� @           |�����>��� � @           |�����>�������� @           ������������ ���� �          ���������|����> @           |�����>��� � @           |�����>�������� @           |�����>���?��?�@           |����>��������� @       �  |����>���?�� @           |����>��������� @           p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ������������?�����?��          ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           ���������|����> @           ��������� @  @           |����>��������� @           |����>���?�� @           |����>��������� @           ������������?�����?��          ���������|����> @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           |����>���?�� @           |����>��������� @           p ���                     ��?������������������������?����          p ��� ��?������?����          ������������������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ������������������                    ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����