�P  XM' +                                                                                                                                               |    |         |    �    �         �    �    �         �   �   �        �   ��  ��        �  ��  ��       d p  ���  ���       �   ���  ���       �� ��� ���      � � � ���    � ��� ���� �     ���� ���   |       ������� @   l  ��?����� D�   8  ���}�� }�      �8����� }�  �  � `���� ��� D `� ����� ��  8 �� A����� C��    �>|������ ��     ��������� �  ���������� �  �  ���@����� �� �  ���`|���| �� �  |��`<���< �� �  <� ���� � � 0 ���~���~    ~ �  ������   � �   ��^ ���    � �  � ��< ���   � � � � �  � ��   � ` � � x@ � � | �   � � b� �   � �     � I  � >  � w    ~  � &  � Z  � ~    8    � � � � �           <      �      ?�      �   ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��   ��   ��   ��   ~�   ~�   ~�   ~�   ��   ��   ��   ��   ~�   ~�   ~�   ~�   ~�   ~�   ~�   ~�   >�   >�   >�   >�  >�  >�  >�  >�  8�  8�  8�  8�  <�  <�  <�  <�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?�  ?�  ?�  ?�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� � � � � � � � �� �� �� �� �� �� �� �� ��  ��  ��  ��  ���.���.���.���.���~���~���~���~�����������������������������������~���~���~���~                                    ' +                                                               �    �         �   �   �        �   �   �            �   �        �   �   �        �       �   `   �   +?   ?�   �       !��  !��        5�  ?��  �   
@  @�  ��  ?�   @ 0  ���  ���  #    �   ��� ���    �  �����     �������      ��
����  �    ���� ��� ��    �������� ��    ��?����� ��
    � ����� ��    � ����� ��>   �|����� ��   |������� ��  ��������� ��   ��������� ��  ��������� ���  ��� ����� ���   �� x���x �� �   �|  ���  �� �   �   ���  �� �   � � ���  �  �  ��� ���       �  �� ��       �   ��  ��       �    ��  ��       �    � �  � �       p    � |  � |  |         � x  � x  �         � |  � |  �        � @  � |  � <        � � � � �     ������������������������������������' + �������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��   p�   p�   p�   p�   ��   ��   ��   ��   p�   p�   p�   p�   p�   p�   p�   p�    �    �    �    �   �   �   �   �  8�  8�  8�  8�  < �  < �  < �  < �  > �  > �  > �  > �  > �  > �  > �  > �  > �  > �  > �  > �  ? �  ? �  ? �  ? �  ?��  ?��  ?��  ?��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� ��� ��� ��� ���������������������������������������������������������������������������������������������������������~���~���~���~������������������������������������' +                   @      `         `  �    � `  �    � `        ` _   _ `       �`  _�   ^ `   � ��`��    `� � ��`��     `  ` ?��`?��     `0 0 ���`���     `�  ?���`���� �   `0� ��� ���� �    @ ��������     `  ?��� ���� �@      ?������@   ��  ?��������         �������� 8       ���������      �ǐ  ��� ��     ��� ���  ��     ��� ���  ��      ��  ���  ��      �   ���  ��      �   ���  ��     �|  ���  ��     ��  ���  ��    ��� ���  G��     3�� ���  ���     ��� ���  �� �   ��  ���  �� �   ��  ���  �� �   �|  ���  �� �   �   ���  �� �   � � ���  �  �  ��� ���       �  �� ��       �   ��  ��       �    ��  ��       �    � �  � �       `    � |  � |  |         � x  � x  �         � |  � |  �        � @  � |  � <        � � � � �                                         ' + ����������������������������������������������������������������������������~����~����~����~��?�>��?�>��?�>��?�>������������������������� �� �� �� �� � � � �    �    �    �    �    �    �    �    �    �    �    �    �   �   �   �   �   �   �   �   �   �   �   �   �   ~�   ~�   ~�   ~�  ~�  ~�  ~�  ~�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ?��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� ��� ��� ��� ���������������������������������������������������������������������������������������������������������~���~���~���~  ��      ��     ��     ��     �' +                                                                                                                           |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��       ��  �  ��   �   @   �  ��  �  �0  <Dx  ?��  ��      ||  ��  ��  @l  �D�  ��  �   �8 ��� ���   |     �9� ��   �   8 �9� ���   �   8 ��� �}�   |       �ǟ ���  ��   8  ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��      �  ���  ��      �| ���  ��    �� ���  ��   ��� ���  ��   0 �� ���  �� � ? ��_ ���  �� � ? ��_ ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ������������������������������������' + �������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ���������������������������������������������������������������������������������� 
����   
����   ����   ����   ��' +                                                                                                                                               |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��       ��  �  ��   �   @   �  ��  �  �0  <Dx  ?��  ��      ||  ��  ��  @l  �D�  ��  �   �8 ��� ���   |     �9� ��   �   8 �9� ���   �   8 ��� �}�   |       �ǟ ���  ��   8  ��� ���  ��      ��� ���  ��      �� ���  ��    �  ���  ��    � / ���  ��    �|k ���  C��    =�y ���  ��     �� ���  �� �  ��_ ���  �� � ? ��_ ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ������������������������������������' + ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������  ����   ~?�      ��     �     �' +                                                                                                                                               |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��        x  ��  ��       d F  ���  ���       ��  ���  ���       �� � � ���    � ��� ���  �   A �ǿ ���   |   @ ��? ���  @  l� �� ���  D�  9  �( ���  }�   �  �8 ���  }�   � �  ���  ��  D �  ���  ��  8 �  ���  ��    � O ���  ��   0 �|� ���  �    0 ��� ���  �  �7 ��� ���  �  � ? ��_ ���  �� � ? ��_ ���  �� � ? ��_ ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �        @   �                            ' + ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ���������������������������������������������������������������������������������������������������� ~������ ~��' +                                                                                                                                                                  �   �        �   �   �            ?�   ?�        0   ��   ��        �   ?�   ��   �    0   �   ��   �    @   �� ��� �     `�  ?��  ���  �@     ?�� �� @   �� ?�� ��� �        �� ��� �        �� ��� �      �ǿ  ��  ��      �� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��   ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      �� ���� ����� F?����� F?����� ' + ������������������������������������������������������������������������������������������������������������������������������������������������������������������?����?����?����?����������������������������������� ��� ��� ��� ��� ��� ��� ��� ���  ���  ���  ���  ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������    �       �       �             ' +                                                                                                                           �    �         �   �   �        �   �   �            �   �        �   �   �        �       �   `   �   +?   ?�   �       !�   !�         5�  ?��  �   
�  @�  ��  ?�   @ F  ���  ���  #    �   ���  ���      �  �� ���      � ��� ���        �� ���   �      ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��   ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ��� ����� ����  ������  ����� ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� G��� G��� G��� G��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������                                    ' +                                                                                                                           |    |         |    �    �         �   �   �        �   ��  ��        �  ��  ��       ��  �  ��   �       �  ��  �   �   D@  ��  ��   @  p  ��  ��  l0  >D�  ?��  �    8  ��  }�|   |   @   �}�  ���   �   �  ��� �}�   |     ��� ���       8 ��� ���         ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��      �  ���  ��    �| ���  ��    �� ���  ��  0 ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ��   ��   ��   ��    ��  ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������� ���� ���� ���� ���� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������  ?����  ?����  ?����  �����  ��' +                                                                                                                           >    >         >    �   �        �   ��   ��        �   ��  ��        `  ��  ��        �  �   ��   �   `  ��  ��   �   �   �  �   A    ��  ;�X  ;��   P  :��  ��  ���   �  �   ��  ���   �  � r �� ���   �    ��? ���       � ��� ���        �� ���   �      ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��  0 ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      �� �� �� �� ��   �    �� �� ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������� ?��� ?��� ?��� ?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ���������������������������������������������������������������������������������� � ?�  ����         a�����  a��' +                                                                                                                                                                   �   �        �   �   �            �   �           ?�   ?�            �   �       @  ��  ��    
  �  ��  ��         ��  ��     `� ���� ����   � � ��������   �    ��� ����   �    ��� ��� ��    ��� ���  �       ��� ���  ��      ��� ���  ��      �� ���  ��      �  ���  ��     �  ���  ��    �| ���  ��    �� ���  ��  0 ��� ���  ��   0 ��� ���  ��   0 ��� ���  �� � 7 �� ���  �� � ? � � ���  �  � ? ��� ���       �  ��� ���       �   ���  ���       �   ��  ��       �   � �  � �       p   � ~  � ~  | |       � ~  � ~  � >       � �  � �  � �       � �  � �  � �            � �  � �      ������������������������������� ' + �������������������������������������������������������������������������������������������������������������������������������������������������������������������?����?����?����?������������������������������������������������������������������� ��� ��� ��� ���  ���  ���  ���  ���  ~��  ~��  ~��  ~�   ~�   ~�   ~�   ~�   >�   >�   >�   >�   >�   >�   >�   >�   ~�   ~�   ~�   ~�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �� 8 �� 8 �� 8 �� 8 �� |�� |�� |�� |�� ��� ��� ��� ����������������������������������������������������������������������������������  ���    ���    ���    ���    �