�P  (#� G �������������������������������������������������������������������������������������������������������������������������                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             ����������������������������� ����������������������������� �                           ������������������������������ �                            �                            �                           ��                            ����������������������������� ����������������������������� �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                        0  
 �                        0  
 �                        0  ������������������������������ �   `` �  �  8       8  
 �   `` �  �  8       8  
 �   `` �  �  8       8  ������������������������������ �  ��� ����� > ` 8x  
 �  ��� ����� > ` 8x  
 �  ��� ����� > ` 8x  ������������������������������ �  �?�� ���� | ��x  
 �  �?�� ���� | ��p  
 �  �?�� ���� | ��x  �������?����������w����������� �  �?�<?� �ǻ��� �����  
 �  �<8<;� �ǁ��p �����  
 �  �?�<?� �ǻ��� �����  �������?�������~7����?������ �  �?�<� �����������=�p  
 �  �<<8q� ��Ǉ0���8=�p  
 �  �?�<� �����������=�p  ���������������|�����?����� �  �|~|���ρ�ϟp����=��  
 �  �|~p� ���� ���<9�p  
 �  �|~|���ρ�ϟp����=��  ���������������������������� �  �<~�������>>���~}��  
 �  �~��p����8 ?��~q��  
 �  �<~�������>>���~}��  �������������>�����?��������� �  �|s������|���~��p  
 �  �8c����x ?��~��`  
 �  �|s������|���~��p  �������������?�|����������o��� �  �9���������x ���q��  
 �  �9�����<�p ���a�`  
 �  �9���������x ���q��  ������ >� �������|F ���� �   �  @      �   
 �                           
 �  �8������x> �����`  ������x  �����<G ��� �   �	   � $     �   
 �                           
 �  �y�����=�p��ø����  ������p� a����8���� �     (        �  @   
 �                           
 �  �<�����>�q������x�  ������0<`� `���C���� �   `@    � d �( @�  
 �                           
 �  �x�ß�����s�����x�  ����� �8< ?� G��� �00���� �  � 78 �@�  @    
 �                           
 �  �}�����߸8����x��9�  �����`><b?� �ǌG��8 ��� �  �@C�@��s� a�    
 �                           
 �  ���Ý����88s���}����  �������?>?�?0�����>�>0���� �  q���@�π8?��@O1�  
 �                           
 �  q�����π8?8��y��1�  ������~������������? ��� �   ��  ` 00 0� q����  
 �                           
 �   ��  ` 00 0� q����  ����������������������~����� �       �       0   q�� p  
 �                           
 �       �       0   q�� p  ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �     >  �        ��|     ������������������������������ �                           
 �                           
 �       �         �B     ������������������������������ �                           
 �                           
 �       �         �B     ������������������������������ �                           
 �                           
 �     p<�Hy��g���B     ������������������������������ �                           
 �                           
 �     �"�H�+ H� �|     ������������������������������ �                           
 �                           
 �     �"�H�� O���QB     ������������������������������ �                           
 �                           
 �     �"�H"�* H@�1B     ������������������������������ �                           
 �                           
 �     �"�0"�* H� �1B     ������������������������������ �                           
 �                           
 �     p<� y�$G��B     ������������������������������ �                           
 �                           
 �                        ������������������������������ �                           
 �                           
 �         � �              ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �     |        @   ���    ������������������������������ �                           
 �                           
 �     B        @   �     ������������������������������ �                           
 �                           
 �     B        @  "     ������������������������������ �                           
 �                           
 �     B�1����0H�A�
"     ������������������������������ �                           
 �                           
 �     |�J@IS(�QA""     ������������������������������ �                           
 �                           
 �     @�! �IR/�a�A"
"     ������������������������������ �                           
 �                           
 �     @��IR( QA""     ������������������������������ �                           
 �                           
 �     @�JAFR(�I�" �     ������������������������������ �                           
 �                           
 �     @�1��D�' D� ���     ������������������������������ �                           
 �                           
 �                         ������������������������������ �                           
 �                           
 �                         ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ��                            ����������������������������� ����������������������������� �                           ������������������������������ �                            �                            �                           ��                             ����������������������������� ����������������������������� �                           ��                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             �                             �                             ������������������������������                              ������������������������������                              ��������������������������������UAUW����UETUW�        ������������UAUW����UETUW�           ����� ���UAUW����UETUW�        ������������UETUW����UETUW�     T      ����� ���U@ UW����U@ UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                  