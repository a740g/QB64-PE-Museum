�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� �� �@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �     @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ����������� �@�       0            ���x� y��       0            ���x� y��       0            ���x� y��       0            �     @�7�������;<��         ���x � |��7�������;<��         ���x � |��7�������;<��         ���x � |��7�������;<������������� �@����6��l�ٳf�         ���x p ~>����6��l�ٳf�         ���x p ~>����6��l�ٳf�         ���x p ~>����6��l�ٳf�         �     @���������3f��         ���x � ~>���������3f��         ���x � ~>���������3f��         ���x � ~>���������3f������������� �@����3�����3f�`         ���x� |�����3�����3f�`         ���x� |�����3�����3f�`         ���x� |�����3�����3f�`         �     @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ����������� �@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �     @�                        ����� ��                        ����� ��                        ����� ��              ��������� �� �@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������M���4�l���ݜp�����T��M���������M���4�l���ݜp�����T��M���������M���4�l���ݜp�����T��M������?������������������������������������5m��w��]��k��[��[S]�]����������5m��w��]��k��[��[S]�]����������5m��w��]��k��[��[S]�]�������?������������������������������������um�o~|-��ݸ.�o��UW]�]����������um�o~|-��ݸ.�o��UW]�]����������um�o~|-��ݸ.�o��UW]�]�������?������������������������������������umvo}�{�������w��UW]�]����������umvo}�{�������w��UW]�]����������umvo}�{�������w��UW]�]�������?�����������������������������������}umu�u�{�]��k��[��n�]�^}��������}umu�u�{�]��k��[��n�]�^}��������}umu�u�{�]��k��[��n�]�^}������?�����������������������������������}um���|,����p�g��n�a��n���������}um���|,����p�g��n�a��n���������}um���|,����p�g��n�a��n�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������0A{�>����������������������������0A{�>����������������������������0A{�>���������������������?����������������������������������������u���;������������������������������u���;������������������������������u���;�����������������������?����������������������������������������}���;������������������������������}���;������������������������������}���;�����������������������?������������������������������������3�}���[�މ�s�nƺ��٘��q��������3�}���[�މ�s�nƺ��٘��q��������3�}���[�މ�s�nƺ��٘��q�����?�����������������������������������u����0�[�����鮺���uַ[{��������u����0�[�����鮺���uַ[{��������u����0�[�����鮺���uַ[{������?�����������������������������������t
������k�~���7뵺ֺ�}۷[{�����t
������k�~���7뵺ֺ�}۷[{�����t
������k�~���7뵺ֺ�}۷[{���?�����������������������������������u�������s������뵺ֺ�}ݷ[{�����u�������s������뵺ֺ�}ݷ[{�����u�������s������뵺ֺ�}ݷ[{���?�����������������������������������u���u���s�����뻺��u��[{��������u���u���s�����뻺��u��[{��������u���u���s�����뻺��u��[{������?������������������������������������;
���A{���s����Y��|q��������;
���A{���s����Y��|q��������;
���A{���s����Y��|q�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������1�8�mfT��p�?�3>6q�������������1�8�mfT��p�?�3>6q�������������1�8�mfT��p�?�3>6q���������?�����������������������������������u��n��{�Z�]�o����w��ծ���w��������u��n��{�Z�]�o����w��ծ���w��������u��n��{�Z�]�o����w��ծ���w������?�����������������������������������u��`��x3n�]�l.�~��઺��������u��`��x3n�]�l.�~��઺��������u��`��x3n�]�l.�~��઺������?�����������������������������������u��o����v�]�k����}����o�����������u��o����v�]�k����}����o�����������u��o����v�]�k����}����o���������?�����������������������������������u��n��{�Z�]�k����u��ծݺ�w��������u��n��{�Z�]�k����u��ծݺ�w��������u��n��{�Z�]�k����u��ծݺ�w������?�������������������������������������q���mgWa�l0�?�>6qݻ�����������q���mgWa�l0�?�>6qݻ�����������q���mgWa�l0�?�>6qݻ�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������o�������������������������������o�������������������������������o�����������������������������?�����������������������������������_���������{����������������������_���������{����������������������_���������{��������������������?�����������������������������������_���������{������������n����������_���������{������������n����������_���������{������������n��������?�����������������������������������O�7{����8yN?2]��c�S�������������O�7{����8yN?2]��c�S�������������O�7{����8yN?2]��c�S�����������?�����������������������������������_��{���k��{5���u����w�}�����������_��{���k��{5���u����w�}�����������_��{���k��{5���u����w�}���������?�����������������������������������_��{�����{tv�}�����z�����������_��{�����{tv�}�����z�����������_��{�����{tv�}�����z���������?�����������������������������������_��{����u�{u���}�����wn����������_��{����u�{u���}�����wn����������_��{����u�{u���}�����wn��������?�����������������������������������_��{.��ku�{u���u����wﯮ����������_��{.��ku�{u���u����wﯮ����������_��{.��ku�{u���u����wﯮ��������?�����������������������������������_�9|�����}v?:����]��������������_�9|�����}v?:����]��������������_�9|�����}v?:����]������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������?����������������������������������?����������������������������������?�������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������������q�8�����������������������������q�8�����������������������������q�8���������?����������������������������������������޿�����������������{���������������޿�����������������{���������������޿�����������������{��������?����������������������������������������߿�����������������{���������������߿�����������������{���������������߿�����������������{��������?������������������������������������7|q�߿�D�9��?1������n���������7|q�߿�D�9��?1������n���������7|q�߿�D�9��?1������n������?�������������������������������������{��؇�[}u������~��|.�8�鮚��������{��؇�[}u������~��|.�8�鮚��������{��؇�[}u������~��|.�8�鮚����?�������������������������������������{�޿�[at���p�����~���}��������{�޿�[at���p�����~���}��������{�޿�[at���p�����~���}����?�������������������������������������{�޿�[]u���u��n�����~������������{�޿�[]u���u��n�����~������������{�޿�[]u���u��n�����~��������?�������������������������������������{��ܿ�[]u���u��n��{���~묺��������{��ܿ�[]u���u��n��{���~묺��������{��ܿ�[]u���u��n��{���~묺����?������������������������������������9|p�⃿[a�9���p��|q�8�����������9|p�⃿[a�9���p��|q�8�����������9|p�⃿[a�9���p��|q�8��������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������?���������������������������������?���������������������������������?�������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?��������������������������������������������������������n���������������������������������n���������������������������������n����������?������������������������������������8|�v>S�O��>S���scO����S�>�?������8|�v>S�O��>S���scO����S�>�?������8|�v>S�O��>S���scO����S�>�?���?�������������������������������������{}u��u�����w���]7�}���t޻��������{}u��u�����w���]7�}���t޻��������{}u��u�����w���]7�}���t޻����?�������������������������������������}��������6�]w�z���޻��������}��������6�]w�z���޻��������}��������6�]w�z���޻����?�����������������������������������u�~ݭ��}������6��]w�wn��}޺������u�~ݭ��}������6��]w�wn��}޺������u�~ݭ��}������6��]w�wn��}޺����?�����������������������������������u�{]���u�ݭ��w���]wﯮ��u޺������u�{]���u�ݭ��w���]wﯮ��u޺������u�{]���u�ݭ��w���]wﯮ��u޺����?�������������������������������������|��?]��ݵ�]����cw����]���?�������|��?]��ݵ�]����cw����]���?�������|��?]��ݵ�]����cw����]���?���?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������o��������{������������������������o��������{������������������������o��������{����������������������?�����������������������������������o���������{������������������������o���������{������������������������o���������{����������������������?�����������������������������������)������h�my��ʜ|���p�?�����������)������h�my��ʜ|���p�?�����������)������h�my��ʜ|���p�?���������?�����������������������������������f�ڻ�}٫o�{w�Zk���]�o��������������f�ڻ�}٫o�{w�Zk���]�o��������������f�ڻ�}٫o�{w�Zk���]�o������������?�����������������������������������n�ڃ�}۫l3{w�Z�=���l.������������n�ڃ�}۫l3{w�Z�=���l.������������n�ڃ�}۫l3{w�Z�=���l.����������?�����������������������������������n�ڿ�|�k�{w��������k��������������n�ڿ�|�k�{w��������k��������������n�ڿ�|�k�{w��������k������������?�����������������������������������n�ڻ�{�k��w�Z뽺�]�k��������������n�ڻ�{�k��w�Z뽺�]�k��������������n�ڻ�{�k��w�Z뽺�]�k������������?����������������������������������������{�l-}����~���l0�7����������������{�l-}����~���l0�7����������������{�l-}����~���l0�7���������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        