�P  `"� M ����������������������������                                                      ���������������������������������������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������                       ���                       ���                           �����������������������������                       ���                       ���                           ��                       ���������������������������������������������������������                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������    P  � @        '����    P  � @        '���      P  � @           �����������������������������    !@  � �        '����    !@  � �        '���      !@  � �           �����������������������������     @   � �        '����     @   � �        '���       @   � �           �����������������������������     S�C�`���g,q�    '����     S�C�`���g,q�    '���       S�C�`���g,q�       �����������������������������     TT �Q@�"�H��     '����     TT �Q@�"�H��     '���       TT �Q@�"�H��        �����������������������������     T �Q@�>�O���    '����     T �Q@�>�O���    '���       T �Q@�>�O���       �����������������������������                      '����                      '���       T �Q@� �H"�        �����������������������������                      '����                      '���      !TR �S@�"�H��        �����������������������������                      '����                      '���      S� ��@��G"q�       �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ����  ���������������������� ���                 '����                      '���   ���                    ����������������������������� ���                 '���� ���                 '���   ��� p �                ����  ����������������������                    '����                    '���   ��� � �                ����  ����������������������                    '����                    '���   ���  �                ����  ����������������������                    '����                    '���   ��� <�I��             ����  ����������������������                    '����                    '���   ��� "�J)              ����  ����������������������                    '����                    '���   ���  "�K�             ����  ����������������������                    '����                    '���   ��� @"�J@             ����  ����������������������                    '����                    '���   ��� �"�2)              ����  ����������������������                    '����                    '���   ��� �<�!��             ����  ����������������������                    '����                    '���   ���                    ����  ���������������������� ���                 '���� ���                 '���         �               ����  ���������������������� ���                 '����                      '���   ���                    �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ����  ���������������������� ���                 '����                      '���   ���                    ����������������������������� ���                 '���� ���                 '���   ���              �    ����  ����������������������                    '����                    '���   ��� �   @       @    ����  ����������������������                    '����                    '���   ���     @       @    ����  ����������������������                    '����                    '���   ���  �q'0O'��,�@    ����  ����������������������                    '����                    '���   ���  �	(�H�����)@    ����  ����������������������                    '����                    '���   ���  �y/�H��"��)�@    ����  ����������������������                    '����                    '���   ���  ��( H��"��)@    ����  ����������������������                    '����                    '���   ���  ��ȠH�����i@    ����  ����������������������                    '����                    '���   ���  �x� O'����@    ����  ����������������������                    '����                    '���   ���  � � H    �  @    ����  ���������������������� ���                 '���� ���                 '���       �  ( 0   �  �    ����  ���������������������� ���                 '����                      '���   ���                    �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ��                       ���������������������������������������������������������                           �����������������������������                       ���                       ���                           �����������������������������                       ���                       ���                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                                                       ��������������������������������������������������������                                          (�(                            ( �� Q8Q��@�Or'�@���D�E� ������������������������������ �(                            (�(                          