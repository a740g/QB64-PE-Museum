�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������}���������_���������������������}���������_���������������������}���������_�����������?�������������������������������������������}w�������������������������������}w�������������������������������}w���������������������?������������������������������������������׻w������������������������������׻w������������������������������׻w���������������������?�����������������������������������S�c<�ݜ��w����MٞS3�N��i������S�c<�ݜ��w����MٞS3�N��i������S�c<�ݜ��w����MٞS3�N��i����?�����������������������������������M�]}��k����u��뽵־���5�[_�������M�]}��k����u��뽵־���5�[_�������M�]}��k����u��뽵־���5�[_�����?�����������������������������������]�A}�ݸ?��w���뽵۾�w�u�]�.������]�A}�ݸ?��w���뽵۾�w�u�]�.������]�A}�ݸ?��w���뽵۾�w�u�]�.����?�����������������������������������]�_}������w��뽵ݾ׷�u��ۮ������]�_}������w��뽵ݾ׷�u��ۮ������]�_}������w��뽵ݾ׷�u��ۮ����?�����������������������������������]�]}��k�}}w�u���=������u�[[�������]�]}��k�}}w�u���=������u�[[�������]�]}��k�}}w�u���=������u�[[�����?�����������������������������������]�c~��}}}��w���Y��;�v��.������]�c~��}}}��w���Y��;�v��.������]�c~��}}}��w���Y��;�v��.����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������~�������������������������������~�������������������������������~�������������?��������������������������������������������������~�������������������������������~�������������������������������~��������������?��������������������������������������������������~�������������������������������~�������������������������������~��������������?�����������������������������������N6�S�q���c�%�˦8~�c"q�4�>�l?������N6�S�q���c�%�˦8~�c"q�4�>�l?������N6�S�q���c�%�˦8~�c"q�4�>�l?����?�����������������������������������5���u�������m�[��~��m���z�k��������5���u�������m�[��~��m���z�k��������5���u�������m�[��~��m���z�k������?�����������������������������������u�^��������m�۬~��m���{~�+�������u�^��������m�۬~��m���{~�+�������u�^��������m�۬~��m���{~�+�����?�����������������������������������u�^�o�����m�ۭ�~��m���{���������u�^�o�����m�ۭ�~��m���{���������u�^�o�����m�ۭ�~��m���{�������?�����������������������������������u۾�u�������m�[-�~��m���z�뫿������u۾�u�������m�[-�~��m���z�뫿������u۾�u�������m�[-�~��m���z�뫿����?�����������������������������������v;�]�q������X�8^��m��7{>�l?������v;�]�q������X�8^��m��7{>�l?������v;�]�q������X�8^��m��7{>�l?����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������_��������������������������������_��������������������������������_������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������S���p�|d�o�N>S3��f8c3����q��������S���p�|d�o�N>S3��f8c3����q��������S���p�|d�o�N>S3��f8c3����q������?�����������������������������������M���[�����o�5������]m溻ٮ��������M���[�����o�5������]m溻ٮ��������M���[�����o�5������]m溻ٮ������?�����������������������������������]��X.��-�o�t�w��Aw۠��������]��X.��-�o�t�w��Aw۠��������]��X.��-�o�t�w��Aw۠������?�����������������������������������]��[����o�u�׷���_{ۯ��������]��[����o�u�׷���_{ۯ��������]��[����o�u�׷���_{ۯ������?�����������������������������������]��[�������u������]mۮ��������]��[�������u������]mۮ��������]��[�������u������]mۮ������?�����������������������������������]��lp��-û�v>�;��8cs������������]��lp��-û�v>�;��8cs������������]��lp��-û�v>�;��8cs����������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������?������������������������������������u�������������������7{����������u�������������������7{����������u�������������������7{�������?������������������������������������}�������������������7{����������}�������������������7{����������}�������������������7{�������?������������������������������������}��c]�~3�q����'�N>�m>�zq���������}��c]�~3�q����'�N>�m>�zq���������}��c]�~3�q����'�N>�m>�zq������?���������������������������������������}]u��ٮ��������5�k�~���������������}]u��ٮ��������5�k�~���������������}]u��ٮ��������5�k�~���������?����������������������������������������]��۠�������t�3}�{��������������]��۠�������t�3}�{��������������]��۠�������t�3}�{�������?����������������������������������������]}�ۯ�������u���|{��������������]}�ۯ�������u���|{��������������]}�ۯ�������u���|{�������?�����������������������������������}u���Yu��ۮ�������u���{���������}u���Yu��ۮ�������u���{���������}u���Yu��ۮ�������u���{�������?�����������������������������������}���e�~7��������v>�m������������}���e�~7��������v>�m������������}���e�~7��������v>�m����������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������7�������������������������������7�������������������������������7����������������������?�����������������������������������o������z�������������������������o������z�������������������������o������z�����������������������?�����������������������������������o������z�������������������������o������z�������������������������o������z�����������������������?�����������������������������������)�Í���z����i�6�c]�}O�a��c��������)�Í���z����i�6�c]�}O�a��c��������)�Í���z����i�6�c]�}O�a��c������?�����������������������������������f���u�{�;�[��v�}]u�7��u��m��������f���u�{�;�[��v�}]u�7��u��m��������f���u�{�;�[��v�}]u�7��u��m������?�����������������������������������n�݅�{z���X.�v��]�w����m��������n�݅�{z���X.�v��]�w����m��������n�݅�{z���X.�v��]�w����m������?�����������������������������������n��u}��z���[��v��]}w��}��m��������n��u}��z���[��v��]}w��}��m��������n��u}��z���[��v��]}w��}��m������?�����������������������������������n��uu�{z���[��y��Yu�w��u��m��������n��uu�{z���[��y��Yu�w��u��m��������n��uu�{z���[��y��Yu�w��u��m������?�������������������������������������Å���{;�lnͻ��e�}w����m����������Å���{;�lnͻ��e�}w����m����������Å���{;�lnͻ��e�}w����m������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������A�/���� ��}������������������������A�/���� ��}������������������������A�/���� ��}��������������?�������������������������������������������_���������}�o����������������������_���������}�o����������������������_���������}�o������������?�������������������������������������������_���������}�o����������������������_���������}�o����������������������_���������}�o������������?��������������������������������������鏻�C��bq�x}��a�)��tL8ό����������鏻�C��bq�x}��a�)��tL8ό����������鏻�C��bq�x}��a�)��tL8ό�����?���������������������������������������w�ۿ]�k������]]of��u��_u�����������w�ۿ]�k������]]of��u��_u�����������w�ۿ]�k������]]of��u��_u�����?����������������������������������������ۿ}��-�����]]�n��u��_u������������ۿ}��-�����]]�n��u��_u������������ۿ}��-�����]]�n��u��_u�����?�����������������������������������u����ۿ}������]]�n��u���u�������u����ۿ}������]]�n��u���u�������u����ۿ}������]]�n��u���u�����?�����������������������������������u���w�ۿ]�뭮����]]on��e��_u�������u���w�ۿ]�뭮����]]on��e��_u�������u���w�ۿ]�뭮����]]on��e��_u�����?������������������������������������և-���cx,m��|w�ca���ݕ�8ߍ��������և-���cx,m��|w�ca���ݕ�8ߍ��������և-���cx,m��|w�ca���ݕ�8ߍ�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������������7���������������������������������7���������������������������������7�������������?�������������������������������������������������c�������������������������������c�������������������������������c���������������?�������������������������������������������������{�������������������������������{�������������������������������{���������������?�����������������������������������&18���N>c1�q��i�{�����������������&18���N>c1�q��i�{�����������������&18���N>c1�q��i�{���������������?�����������������������������������o��[�{5��~���릺�{�;���������������o��[�{5��~���릺�{�;���������������o��[�{5��~���릺�{�;�������������?�����������������������������������n�o�{t�p���.�zu����������������n�o�{t�p���.�zu����������������n�o�{t�p���.�zu��������������?�����������������������������������m����{u��n�o����{�����������������m����{u��n�o����{�����������������m����{u��n�o����{���������������?�����������������������������������m��[�{u��n���ˮ��{�����������������m��[�{u��n���ˮ��{�����������������m��[�{u��n���ˮ��{���������������?�����������������������������������n���}v?c��q�,n�{�:���������������n���}v?c��q�,n�{�:���������������n���}v?c��q�,n�{�:�������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        