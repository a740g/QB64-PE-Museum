�P  @u ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                               ��                               ��                               ��                               ��                               ��                               ��                               ��              ����������������@��                           ���                           ���                           ���                           @��                            s���                            s���                            s���           ����������������@��                            y���                            y���                            y���                            @����y�                         |�����y�                         |�����y�                         |�����y�        ����������������@�gm��                         ~>�gm��                         ~>�gm��                         ~>�gm��                         @�fm�|�                         ~>�fm�|�                         ~>�fm�|�                         ~>�fm�|�        ����������������@��m���                         |���m���                         |���m���                         |���m���                         @�6m�Ͱ                         y��6m�Ͱ                         y��6m�Ͱ                         y��6m�Ͱ        ����������������@�6m�}�                         s��6m�}�                         s��6m�}�                         s��6m�}�                         @�                               ��                               ��                               ��              ����������������@�                               ��                               ��                               ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ���� ��������������������������������� ��������������������������������� ������������������������������                               ����������������������������������������������������������������������������������������������������������  ��                            �������������������������������������������������������������������������������������������������������  ?��                            ��������w����������������������������������w����������������������������������w���������������������������  ��                            ��������w����������������������������������w����������������������������������w���������������������������  ��                            ��������t��Li���1���ӎ|8�O���������������t��Li���1���ӎ|8�O���������������t��Li���1���ӎ|8�O��������  ��                            ��������s]�ۦ�޻뮻ڻ����]7���������������s]�ۦ�޻뮻ڻ����]7���������������s]�ۦ�޻뮻ڻ����]7��������  ��                            ��������wA��.�޻��ڃ݆��Aw���������������wA��.�޻��ڃ݆��Aw���������������wA��.�޻��ڃ݆��Aw��������  ��                            ��������w_���޺믻ڿ�w}��w���������������w_���޺믻ڿ�w}��w���������������w_���޺믻ڿ�w}��w��������  ��                            ��������w]�ۮ�>�뮻ڻ�u��]w���������������w]�ۮ�>�뮻ڻ�u��]w���������������w]�ۮ�>�뮻ڻ�u��]w��������  ��                            ��������wc���n�~�1���݆|8�w���������������wc���n�~�1���݆|8�w���������������wc���n�~�1���݆|8�w��������  ��                            �������������������������������������������������������������������������������������������������������  ��                            ����������������������������������������������������������������������������������������������������������  ��                            ����������������������������������������������������������������������������������������������������������  ��                            ����������������������������������������������������������������������������������������������������������  ��                            ������������������~���������������������������������~���������������������������������~����������������  ��                            �������������������������������������������������������������������������������������������������������  ��                            ����������������������������������������������������������������������������������������������������  ��                            ��������4�c��c���mf�1���~4�N��������������4�c��c���mf�1���~4�N��������������4�c��c���mf�1���~4�N�������  ��                            ��������պ�w�]���mZon����}5�[�������������պ�w�]���mZon����}5�[�������������պ�w�]���mZon����}5�[������  ��                            ����������w�]���Un�n��X=�au�o���������������w�]���Un�n��X=�au�o���������������w�]���Un�n��X=�au�o������  ��                            ��������վ�w�]���Uv�n��[��]u���������������վ�w�]���Uv�n��[��]u���������������վ�w�]���Uv�n��[��]u��������  ��                            ��������պ�w����ϻZ�n�����]u�[�������������պ�w����ϻZ�n�����]u�[�������������պ�w����ϻZ�n�����]u�[������  ��                            ��������������/�f��ü~7av�������������������/�f��ü~7av�������������������/�f��ü~7av������  /��                            ���� ��������������������������������� ��������������������������������� ������������������������������                                ���� ����������������������?���������� ����������������������?���������� ����������������������?�������  ��                            ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ���        �        �        ������        �        �        ������        �        �        ����                                 �������������������������������������������������������������������������������������������������  �������� �������� ��������  �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         ����������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �����������������������N8�����������������������������N8�����������������������������N8�������  @        @        @         �������o���������������5�_������������o���������������5�_������������o���������������5�_������  @        @        @         ���������������W�������u�_��������������������W�������u�_��������������������W�������u�_������  @        @        @         �����������������������u������������������������������u������������������������������u��������  @        @        @         �������o��������������]u�_������������o��������������]u�_������������o��������������]u�_������  @        @        @         �����������������������v8�����������������������������v8�����������������������������v8�������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         �������������������������������������������������������������������������������������������������  @        @        @         ���        �        �        ������        �        �        ������        �        �        ����  �������� �������� ��������  ���        �        �        ������        �        �        ������        �        �        ����                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                