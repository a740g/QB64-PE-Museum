�3  �x ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �           �<  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ���������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��          ��  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��@         
��  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��            ��_�                                                        �����            ��_�                                                        �����            ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �       ��_�                                                        �����     �       ��_�                                                        �����     �       ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �       ��_�                                                        �����     �       ��_�                                                        �����     �       ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �       ��_�                                                        �����     �       ��_�                                                        �����     �       ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �y͠    ��_�                                                        �����     �y͠    ��_�                                                        �����     �y͠    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �}�    ��_�                                                        �����     �}�    ��_�                                                        �����     �}�    ��_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �}�   ���_�                                                        ������   �}�   ���_�                                                        ������   �}�   ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �}�   ���_�                                                        ������   �}�   ���_�                                                        ������   �}�   ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �T"    ���_�                                                        ������   �T"    ���_�                                                        ������   �T"    ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �T�    ���_�                                                        ������   �T�    ���_�                                                        ������   �T�    ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���   �U"    ���_�                                                        ������   �U"    ���_�                                                        ������   �U"    ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ��     �U�    ��_�                                                        �����     �U�    ��_�                                                        �����     �U�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �U�    ��_�                                                        �����     �U�    ��_�                                                        �����     �U�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �U�    ��_�                                                        �����     �U�    ��_�                                                        �����     �U�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��     �T�    ��_�                                                        �����     �T�    ��_�                                                        �����     �T�    ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ���           ���_�                                                        ������           ���_�                                                        ������           ���_�                                                        ��� �_�����������<  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                                                        �����              ��_�                                                        �����              ��_�                                                        ��� ��_������������  �������������������������������������������������������π! ��              ��_�                   �               >                  �����              ��_�                   �               >                  �����              ��_�                   �               >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                   �               >                  �����              ��_�                   �               >                  �����              ��_�                   �               >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                   �               >                  �����              ��_�                   �               >                  �����              ��_�                   �               >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                   �               >                  �����              ��_�                   �               >                  �����              ��_�                   �               >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                   �               >                  �����              ��_�                   �               >                  �����              ��_�                   �               >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                  ���              >                  �����              ��_�                  ���              >                  �����              ��_�                  ���              >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                  ���              >                  �����              ��_�                  ���              >                  �����              ��_�                  ���              >                  ��� ��_������������  �������������������������������������������������������π! ��              ��_�                  ���              >                  �����              ��_�                  ���              >                  �����              ��_�                  ���              >                  ��� �@         
�<  �������������������������������������������������������π! ���           ���_�                  ���              >                  ������           ���_�                  ���              >                  ������           ���_�                  ���              >                  ��� ������������<  �������������������������������������������������������π! ���           ���_�                  ���              >                  ������           ���_�                  ���              >                  ������           ���_�                  ���              >                  ��� �          �<  �������������������������������������������������������π! ���           ���_�                  ���               >                  ������           ���_�                  ���               >                  ������           ���_�                  ���               >                  ��� �������������<  �������������������������������������������������������π! ���           ���_�                  ���               >                  ������           ���_�                  ���               >                  ������           ���_�                  ���               >                  ��� �           �<  �������������������������������������������������������π! ���           ���_�                  ���               >                  ������           ���_�                  ���               >                  ������           ���_�                  ���               >                  ��� �������������<  �������������������������������������������������������π! ��              ��_�                  ���               >                  �����              ��_�                  ���               >                  �����              ��_�                  ���               >                  ��� ���������������  �������������������������������������������������������π! �������������������_�                  ���               >                  ����������������������_�                  ���               >                  ����������������������_�                  ���               >                  ���?�������������������������������������������������������������������������π! �������������������_�                  ���               >                  ����������������������_�                  ���               >                  ����������������������_�                  ���               >                  ���                  �������������������������������������������������������π! ����           ���_�                  ���               >                  �������           ���_�                  ���               >                  �������           ���_�                  ���               >                  ���               @  �������������������������������������������������������π! ����           ���_�                  ���               >                  �������           ���_�                  ���               >                  �������           ���_�                  ���               >                  ���               @  �������������������������������������������������������π! ���           ���_�                  ���               >                  ������           ���_�                  ���               >                  ������           ���_�                  ���               >                  ���              �  �������������������������������������������������������π! ����           ��z_�                  ���               >                  �������           ��z_�                  ���               >                  �������           ��z_�                  ���               >                  ��� � ������������ �������������������������������������������������������π! ����           ��_�                  � �?���������>                  �������           ��_�                  � �?���������>                  �������           ��_�                  � �?���������>                  ���!�           � ��������������������������������������������������������π! ����           ��_�                  � �?���������>                  �������           ��_�                  � �?���������>                  �������           ��_�                  � �?���������>                  ���!� ����������� ��������������������������������������������������������π! �w��           ��_�                  � �?���������>                  ����w��           ��_�                  � �?���������>                  ����w��           ��_�                  � �?���������>                  ���!p @         
� ��������������������������������������������������������π! ����           ��z_�                  � �?���������>                  �������           ��z_�                  � �?���������>                  �������           ��z_�                  � �?���������>                  ��� � _����������� �������������������������������������������������������π! ���           ���_�                  � �?���������>                  ������           ���_�                  � �?���������>                  ������           ���_�                  � �?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  �������           ���_�                  � �?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  �������           ���_�                  ���?���������>                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���> |��|  > � >                  �������           ���_�                  ���> |��|  > � >                  �������           ���_�                  ���> |��|  > � >                  ���   _�����������  �������������������������������������������������������π! ����           ���_�                  ���> |��|  > � >                  �������           ���_�                  ���> |��|  > � >                  �������           ���_�                  ���> |��|  > � >                  ���   _�����������  �������������������������������������������������������π! ����         ���_�                  ���> |��|  > � >                  �������         ���_�                  ���> |��|  > � >                  �������         ���_�                  ���> |��|  > � >                  ���   _�����������  �������������������������������������������������������π! ����   �      ���_�                  ���> |��|  > � >                  �������   �      ���_�                  ���> |��|  > � >                  �������   �      ���_�                  ���> |��|  > � >                  ���   _�����������  �������������������������������������������������������π! ����   �      p  :_�                  ���> |��|  > � >                  �������   �      p  :_�                  ���> |��|  > � >                  �������   �      p  :_�                  ���> |��|  > � >                  ���   _�����������  $�������������������������������������������������������π! ����   �      p  :_�                  � �> |��| �� � >                  �������   �      p  :_�                  � �> |��| �� � >                  �������   �      p  :_�                  � �> |��| �� � >                  ���   _���������������������������������������������������������������������π! ����   �y͠   p  :_�                  � �> |��| �� � >                  �������   �y͠   p  :_�                  � �> |��| �� � >                  �������   �y͠   p  :_�                  � �> |��| �� � >                  ���   _���������������������������������������������������������������������π! ����   �}�   pp:_�                  � �> |��| �� � >                  �������   �}�   pp:_�                  � �> |��| �� � >                  �������   �}�   pp:_�                  � �> |��| �� � >                  ���   _���������������������������������������������������������������������π! ����   �}�   p"�:_�                  � �> |��| �� � >                  �������   �}�   p"�:_�                  � �> |��| �� � >                  �������   �}�   p"�:_�                  � �> |��| �� � >                  ���   _���������������������������������������������������������������������π! ����   �}�   p"�:_�                  � �> |��| �� � >                  �������   �}�   p"�:_�                  � �> |��| �� � >                  �������   �}�   p"�:_�                  � �> |��| �� � >                  ���   _���������������������������������������������������������������������π! ����   �T"    p"�:_�                  � �> |��| > � >                  �������   �T"    p"�:_�                  � �> |��| > � >                  �������   �T"    p"�:_�                  � �> |��| > � >                  ���   _���������������������������������������������������������������������π! ����   �T�    p"�:_�                  � �> |��| > � >                  �������   �T�    p"�:_�                  � �> |��| > � >                  �������   �T�    p"�:_�                  � �> |��| > � >                  ���   _���������������������������������������������������������������������π! ����   �U"    p"�:_�                  � �> |��| > � >                  �������   �U"    p"�:_�                  � �> |��| > � >                  �������   �U"    p"�:_�                  � �> |��| > � >                  ���   _���������������������������������������������������������������������π! ����   �U�   p"�:_�                  � �> |��| > � >                  �������   �U�   p"�:_�                  � �> |��| > � >                  �������   �U�   p"�:_�                  � �> |��| > � >                  ���   _���������������������������������������������������������������������π! ����   �U�   p"�:_�                  � �> |��| > � >                  �������   �U�   p"�:_�                  � �> |��| > � >                  �������   �U�   p"�:_�                  � �> |��| > � >                  ���   _���������������������������������������������������������������������π! ����   �U�   pp:_�                  � �> |��|����                   �������   �U�   pp:_�                  � �> |��|����                   �������   �U�   pp:_�                  � �> |��|����                   ���   _���������������������������������������������������������������������π! ����   �T�   p  :_�                  � �> |��|����                   �������   �T�   p  :_�                  � �> |��|����                   �������   �T�   p  :_�                  � �> |��|����                   ���   _���������������������������������������������������������������������π! ����           p  :_�                  � �> |��|����                   �������           p  :_�                  � �> |��|����                   �������           p  :_�                  � �> |��|����                   ���   _���������������������������������������������������������������������π! ����           p  :_�                  � �> |��|����                   �������           p  :_�                  � �> |��|����                   �������           p  :_�                  � �> |��|����                   ���   _���������������������������������������������������������������������π! ����           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   ���   _���������������������������������������������������������������������π! ����           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   ���   _�����������  �������������������������������������������������������π! ����           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   �������           ���_�                  � �> |��|����                   ���   _�����������  �������������������������������������������������������π!   �C������ ������������ ���               ���������� ������������            /I�  �
�  ж?���-�;� ������������ /I�  �
�      �w� ������H�Q� ������������     ��w�             ���������� ������������     �              ���������� ������������     �                ���������� ������������     �              ���������� ������������     �              ���������� ������������     �              ���������� ���������������������          ���������� ����������������������          ���������� ����������������������          ���������� ����������������������          ?���������� ����������������������            ?���������� ����������������������      >      ����������������������@����������      ��     ������������          @                 x?�����?������������          @                 �         ��     ����� �����                                    ������������                    