�P�`;c ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                               ��                               ��                               ��                               ��                               ��                               ��                               ��              ����������������@��                             ���                             ���                             ���                             @�`                             s��`                             s��`                             s��`            ����������������@�`                             y��`                             y��`                             y��`                             @�o�>                           |��o�>                           |��o�>                           |��o�>          ����������������@�lٻ                           ~>�lٻ                           ~>�lٻ                           ~>�lٻ                           @�l߳                           ~>�l߳                           ~>�l߳                           ~>�l߳          ����������������@�l�3                           |��l�3                           |��l�3                           |��l�3                           @�lٳ                           y��lٳ                           y��lٳ                           y��lٳ          ����������������@�Ϗ3                           s��Ϗ3                           s��Ϗ3                           s��Ϗ3                           @�                              ��                              ��                              ��             ����������������@�                              ��                              ��                              ��                              @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                ��                                ��                                ��                                 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                ��                                ��                                ��                                 �����������������������������������������������������������������������������������������������������������                                 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������           ~����������������������           ~����������������������           ~�                                 ���������������������������������~���������������������������������~���������������������������������~�                    �������������������������������������������~��������������������������������~��������������������������������~�                         @    ���������������������������������~���������������������������������~���������������������������������~�                         @    ���������������������������������~���������������������������������~���������������������������������~�                         @    ������s�n�����ӌ���������������~������s�n�����ӌ���������������~������s�n�����ӌ���������������~�                         @    ��5w��k���]��M���u�������������~��5w��k���]��M���u�������������~��5w��k���]��M���u�������������~�                         @    ����h7���A��݅���������������~����h7���A��݅���������������~����h7���A��݅���������������~�                         @    �����k����_���u��}���?��������~�����k����_���u��}���?��������~�����k����_���u��}���?��������~�                         @    ���w��k���]��]u��u���������޷��~���w��k���]��]u��u���������޷��~���w��k���]��]u��u���������޷��~�                         @    �����ls������݅�����������ޯ��~�����ls������݅�����������ޯ��~�����ls������݅�����������ޯ��~�                         @    ������������������������ӎ7��ޟ��~������������������������ӎ7��ޟ��~������������������������ӎ7��ޟ��~�                         @    ������������������������Mu���ޟ��~������������������������Mu���ޟ��~������������������������Mu���ޟ��~�                         @    ������������������������]|��ޯ��~������������������������]|��ޯ��~������������������������]|��ޯ��~�                         @    ������������������������]}���޷��~������������������������]}���޷��~������������������������]}���޷��~�                         @    ������������������������]u���޻��~������������������������]u���޻��~������������������������]u���޻��~�                         @    ��3��?����ާ�1��q����8]�7�����~��3��?����ާ�1��q����8]�7�����~��3��?����ާ�1��q����8]�7�����~�                         @    ����Z����m�ޚ���{��������������~����Z����m�ޚ���{��������������~����Z����m�ޚ���{��������������~�                         @    ����o���m�޺���{��������������~����o���m�޺���{��������������~����o���m�޺���{��������������~�                         @    ���������mv޺���{��������������~���������mv޺���{��������������~���������mv޺���{��������������~�                         @    ����Z����mw>��ˮ�{��������������~����Z����mw>��ˮ�{��������������~����Z����mw>��ˮ�{��������������~�                         @    ��7��7��/m�~�,1�xp�_������������~��7��7��/m�~�,1�xp�_������������~��7��7��/m�~�,1�xp�_������������~�                         @    ��������������������������������~��������������������������������~��������������������������������~�                         @    ���������������������������������~���������������������������������~���������������������������������~�                         @    ����������������������           ~����������������������           ~����������������������           ~�                    ���������������������������������           ~����������������������           ~����������������������           ~�                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          ���������������������������������������������������������������������������������������������������������������������������������������������                              -                          x     x     x     x     �     �     �     �     �     �     �     �     ��3�  ��3�  ��3�  ��3�  x6`  x6`  x6`  x6`  ���  ���  ���  ���  ��   ��   ��   ��   ͘�`  ͘�`  ͘�`  ͘�`  x���  x���  x���  x���                                                  ��������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ������������������������������������-                          x   0 x   0 x   0 x   0 �   0 �   0 �   0 �   0 �   x �   x �   x �   x ��3�xp��3�xp��3�xp��3�xpx6`��x6`��x6`��x6`������`����`����`����`�� �0�� �0�� �0�� �0͘�a��͘�a��͘�a��͘�a��x����px����px����px����p                                                ����������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������