�P  �>  P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � @H                      �{���������������                     B�! ��P�a��                     B� ��^�y���                    ��n���߀���������                    �K����߀���������                     K�����������0�                    �{����߀���������                    ��q�������������                    O������B�!B0�  �{���            �������?����������                    ������������������            �{���  O������B�!B�                    O������O������                    ������������������               �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P - ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        �        �        �        ��9�{��-���9�{��-���9�{��-���9�{��-���9�	��$��9�	��$��9�	��$��9�	��$�        �        �        �        �        �        �        �        ��0    ���0    ���0    ���0    ��        �        �        �        �        �        �        �        ���    ����    ����    ����    ��        �        �        �        �        �        �        �        ���    ����    ����    ����    ����    ����    ����    ����    ��        �        �        �        �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P ���������������������������                    ������������������                    ������������������                    ������������������                    ������������������                    ���������          ���������          ������������������          ������������������                              ������������������          ������������?���                     8p 8  Ǐ�������Ǐ�������          ������������������                     �� G� #� p;�����p;�����          �?�����~���g���~    �           � P)(��
@}�����`�}��׃`�       � �'����	�{o�}����    7�           � "��AD�z���w����z }w��� ^  � @;�#�����v���w����    w�      @  ;�
!E��Pu������ �t  ���]  .  @  �{�P���������t  �  }  >             @     
!E��Pu������{��t  ���]  .  @  �  P~!���~u������{��    ��      @  �  P
!E��Pu������{��t  ���]  .  @  �  P~!���~u������{��    ��      @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P��E������u��������t  �  ]  .��@��������������w���������             @     x  |  >  ������������������x  |  >  ������������������                              ������������������          ������������������                    x  |  >  ������������������          ���������w���������             @     ��E������t  �  }  >t  �  ]  .   @     ~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P��E������t  �  }  >t  �  ]  .   @     ~!���~u������{��            @  �  P
!E����u������{��t  �  ]{��  @  �  P~!�����u������{��       {��  @  �  P
!E���Pu������{�~t  �  ]{�.  @  � �~!����~u������{�~       {�   @  � �
!E���Pu������{�~t  �  ]{�.  @  � �~!����~u������{�~       {�   @  � ���E������u��������t  �  ]  .��@��������������w���������             @       D  "  w���������w���������   @     ������������������          ���������          ������������������          ������������������                    ���������                              ���������w���������             @       D  "  w���������w���������   @     ���������t  �  }  >             @     
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P���������t  �  }  >             @     
!E��Pu������{�~t  �  ]�.  @  � w�~!���~u������{�~       �   @  � w�
!E��Pu������{�~t  �  ]�.  @  � w�~!���~u������{�~       �   @  � w�
!E��Pu������{�~t  �  ]�.  @  � w�~!���~u������{�~       �   @  � w�
!E��Pu������{�~t  �  ]�.  @  � w����������u��������          ��@�����  D  "  w���������w���������   @     ���������w���������             @     x  |  >  ������������������x  |  >  ������������������                              ������������������          ������������������                    x  |  >  ������������������          ���������w���������             @     ��E������t  �  }  >t  �  ]  .   @     �'����~u������{��� �       @  �  P�'E���Pu������{��u��� ]  .  @  �  P�'����~u������{��� �       @  �  P��E���Pu������{��u�޺� ]  .  @  �  P������~u������{���� �       @  �  P��E���Pu������{��u�޺� ]  .  @  �  P������~u������{���� �       @  �  P��E������t  �  }  >t  �  ]  .   @     ������~u������{���� �       @  �  P��E���Pu������{��u�޺� ]  .  @  �  P�����~u������{����         @  �  P��E��Pu������{��u�޺  ]  .  @  �  P~����~u������{�� �         @  �  P
�E��Pu������{��t޺  ]  .  @  �  P~����~u������{�� �         @  �  P��E������u��������t  �  ]  .��@��������������w���������             @       D  "  w���������w���������   @     ������������������          ���������          ������������������          ������������������                    ���������                              ���������w���������             @       D  "  w���������w���������   @     ���������t  �  }  >             @     
!E��Pu�����{��t  � o]{�. �@  �  P~!���~u�����{��     o {�  �@  �  P
!E��Pu�����{��t  � o]{�. �@  �  P~!���~u�����{��     o {�  �@  �  P
!E��Pu�����{��t  � o]{�. �@  �  P~!���~u�����{��       {�  �@  �  P
!E��Pu�����{��t  �  ]{�. �@  �  P���������t  �  }  >             @     
!E��Pu������{��t  �  ]{�.  @  �  P~!���~u������{��       {�   @  �  P
!E��Pu������{��t  �  ]{�.  @  �  P~!���~u������{��       {�   @  �  P
!E��Pu������{��u� �  ]{�.  @  �  P~!���~u������{���          @  �  P
!E��Pu������{��u� �  ]  .  @  �  P���������u��������          ��@�����  D  "  w���������w���������   @     ���������w���������             @     x  |  >  ������������������x  |  >  ������������������                              ������������������          ������������������                    x  |  >  ������������������          ���������w���������             @     ��E������t  �  }  >t  �  ]  .   @     ~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P��E������t  �  }  >t  �  ]  .   @     ~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{�� �         @  �  P
!E��Pu������{��t޺  ]  .  @  �  P~!���~u������{�� �         @  �  P��E������u��������t  �  ]  .��@��������������w���������             @       D  "  w���������w���������   @     ������������������          ���������          ������������������          ������������������                    ���������                              ���������w���������             @       D  "  w���������w���������   @     ���������t  �  }  >             @     
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E����Pu������{��t  ���]  .  @  �  P~!�����~u������{��    ��      @  �  P
/E����Pu������{��t ���]  .  @  �  P���������t  �  }  >             @     
/E����Pu������{��t ���]  .  @  �  P~/�����~u������{��   ��      @  �  P
/E����Pu������{��t ���]  .  @  �  P�/�����~u������{��� ��      @  �  P�/E����Pu������{��u����]  .  @  �  P�/�����~u������{��� ��      @  �  P�/E����Pu������{��u����]  .  @  �  P���������u��������          ��@�����  D  "  w���������w���������   @     ���������w���������             @     x  |  >  ������������������x  |  >  ������������������                              ������������������          ������������������                    x  |  >  ������������������          ���������w���������             @     ��E������t  �  }  >t  �  ]  .   @     ~!�P��~t������{��    ��   � @  �  P
!EP��Pt������{��t  ���]  � @  �  P~!�P��~t������{��    ��   � @  �  P
!EP��Pt������{��t  ���]  � @  �  P~!�P��~t������{��    ��   � @  �  P
!EP��Pt������{��t  ���]  � @  �  P~!�����~t������{��    ��     @  �  P��E������t  �  }  >t  �  ]  .   @     ~!���~t������{��       {�  @  �  P
!E��Pt������{��t  �  ]{�. @  �  P~!���~u������{��       {�   @  �  P
!E��Pu������{��t  �  ]{�.  @  �  P~!���~u������{��       {�   @  �  P
!E��Pu������{��t  � ]{�.  @  �  P~!���~u������{��   � {�   @  �  P��E������u��������t  �  ]  .��@��������������w���������             @       D  "  w���������w���������   @     ������������������          ���������          ������������������          ������������������                    ���������                              ���������w���������             @       D  "  w���������w���������   @     ���������t  �  }  >             @     
!E��Pu�����{��t ��]@ .  ]@  �  P~!���~u�����{��   �       ]@  �  P
!E��Pu�����{��t  �  ]  .  _@  �  P~!���~u�����{��            _@  �  P
!E��Pu�����{��t  �  ]  .  _@  �  P~!���~u�����{��            _@  �  P
!E��Pu�����{��t  �  ]  .  _@  �  P���������t  �  }  >             @     
!E��Pu�����{��t  �  ]  .  _@  �  P~!�����~u�����{��    ��      _@  �  P
!E��Pu�����{��t  ���]  .  _@  �  P~!�����~u�����{��    ��      _@  �  P
!E��Pu�����{��t  ���]  .  _@  �  P~!�����~u������{��    ��      @  �  P
!E��Pu������{��t  ���]  .  @  �  P���������u��������          ��@�����  D  "  w���������w���������   @     ���������w���������             @     x  |  >  ������������������x  |  >  ������������������                              ������������������          ������������������                    x  |  >  ������������������          ���������w���������             @     ��E������t  �  }  >t  �  ]  .   @     ~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @  �  P
!E��Pu������{��t  �  ]  .  @  �  P~!���~u������{��            @ �  P
!E��Pu������{��t  �  ]  .  @ �  P~!���~u������{��            @ �  P��E������t  �  }  >t  �  ]  .   @     ~!���~u������{��            @ �  P
!E��Pu������{��t  �  ]  .  @ �  P~!���~u������{��            @ �  P
!E��Pu������{��t  �  ]  .  @ �  P~!���~u������{��            @ �  P
!E��Pu������{��t  �  ]  .  @ �  P~!���~u������{��            @ �  P��E������u��������t  �  ]  .��@��������������w���������             @               ������������������          ������������������          ���������          ������������������          ������������������                    ���������                              ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                              ������������������          ������������������                    ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����