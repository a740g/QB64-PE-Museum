�P   AU � ������������������������������������������������������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         �������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ��/����������/����������/���������         ��.����������.����������.���������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         ����������������������������������         ����������������������������������         ���Ɵ���������Ɵ���������Ɵ�������         ����o����������o����������o�������         ����������������������������������         ����������������������������������         ����������������������������������         ��a����������a����������a���������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         ����������������������������������         ���v?���������v?���������v?�������         ���u����������u����������u��������         ��a���������a���������a��������         ��]����������]����������]���������         ��]����������]����������]���������         ����?����������?����������?�������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         ����������������������������������         ���v?�?�������v?�?�������v?�?�����         ���u�v��������u�v��������u�v������         ��a�w������a�w������a�w�����         ��]���������]���������]��������         ��]����������]����������]���������         ����>�?��������>�?��������>�?�����         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �         0�         0�         0����������������������������������������������������������������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         �������������������������������         �������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ��_����������_����������_���������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         �������������������������������         �������������������������������         ����������������������������������         �������������������������������         �������������������������������         �������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         �         0�         0�         0����������������������������������������������������������������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ��~����������~����������~���������         ����������������������������������         ����������������������������������         ��ڟ���������ڟ���������ڟ��������         ��ڿ���������ڿ���������ڿ��������         �������������������������������         �������������������������������         ��ڿ���������ڿ���������ڿ��������         ��Z����������Z����������Z���������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������                                          �����������������  ��     5 9 ��������������������������������������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     �������������������     ����������������������     ����������������������     ����������������������     ����������������������     ��n�����n�����n����     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     �������������������     ����������������������     ����������������������     ���o�����o�����o���     ���o�����o�����o���     ���o�����o�����o���     ���o�����o�����o���     ����������������������     ��q������q������q�����     ����������������������     �������������������     ����������������������     ����������������������     ����������������������     �������������������     ����������������������     ����������������������     ����������������������     ��~������~������~�����     ���݃�����݃�����݃���     �������������������     �������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������     ����������������������                          �������W + ������������������������������������������������������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������         ����������������������������         �������������������������������         ���c���������c���������c�������         ���]u�~�������]u�~�������]u�~�����         ��AA}�����AA}�����AA}����         ��__}�����__}�����__}����         ��]]u�����]]u�����]]u����         ���c��������c��������c������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ��}���������}���������}��������         ����{����������{����������{�������         �������������������������������         ���O�������O�������O�����         ���_~��o������_~��o������_~��o����         ���_~��������_~��������_~������         ���_~���������_~���������_~�������         ���_z��o������_z��o������_z��o����         ��ao�������ao�������ao������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������         ����������������������������������                                          �����������                           ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��������������������������������������������������������b 9 ��������������������������������������������������������������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @��W������������W������������W�����������           @����������������������������������������           @����������������������������������������           @���>�2�4�ko�����>�2�4�ko�����>�2�4�ko���           @�������_�o���������_�o���������_�o���           @��������\+o����������\+o����������\+o���           @��������[�o����������[�o����������[�o���           @�����ֽ�[���������ֽ�[���������ֽ�[�����           @���>�6�7l+������>�6�7l+������>�6�7l+����           @����������������������������������������           @�������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @��W������������W������������W�����������           @�������������������������������������           @����w�����������w�����������w��������           @���?w,q��������?w,q��������?w,q������           @����v�k����������v�k����������v�k�������           @���߮k�������߮k�������߮k�����           @���߮�k������߮�k������߮�k����           @������k�����������k�����������k������           @���?��p��������?��p��������?��p������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @�������������������������������������           @�������������������������������������           @�������������������������������������           @����]��q�������]��q�������]��q����           @�����]w�����������]w�����������]w�������           @����k���������k���������k������           @��/��k��������/��k��������/��k�������           @��.��ww��������.��ww��������.��ww�������           @����w����������w����������w�������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @����������������������������������������           @                                       �������������a 9 ������������ ������������ ������������ ������������������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ���9��e�9���� ��9��e�9���� ��9��e�9���� �           ���ֶ�t����� ��ֶ�t����� ��ֶ�t����� �           ���۶��u����� ��۶��u����� ��۶��u����� �           ���ݶ��u����� ��ݶ��u����� ��ݶ��u����� �           ���ֶ˭u����� ��ֶ˭u����� ��ֶ˭u����� �           �����,u������ ����,u������ ����,u������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ���������+�� ��������+�� ��������+�� �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           �����18��� ����18��� ����18��� �           ���������xj�� ��������xj�� ��������xj�� �           ���݅���{�� ��݅���{�� ��݅���{�� �           ����u����{��� ���u����{��� ���u����{��� �           ����u����{��� ���u����{��� ���u����{��� �           ���c�6���� ��c�6���� ��c�6���� �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ���w�������� ��w�������� ��w�������� �           ���p�t�t�8��� ��p�t�t�8��� ��p�t�t�8��� �           ����]u��V�Z�� ���]u��V�Z�� ���]u��V�Z�� �           ����]u��V�f�� ���]u��V�f�� ���]u��V�f�� �           ���7]u�7V�f�� ��7]u�7V�f�� ��7]u�7V�f�� �           ����]e��V�[�� ���]e��V�[�� ���]e��V�[�� �           �������V�Z�� ������V�Z�� ������V�Z�� �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           ������������� ������������ ������������ �           �                                       �������������    