�P   ˀ� ��������������?�����������������������?��������������                        �    �����@   �������    �����@   ��������                           ?�������     �������     �������     �������     �                           BN     �     �     8          �     �     8     $                        �~�����������p����������������������p��������������                         8   ?������@   #�������   ?������@   #��������                            ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8                             ���������������������������������������������������                        @�   �������@  �8������   �������@  �8�������                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      D                        ��7���������������������g�����������������������g����                        �8@  f �����D  ` ������@  f �����D  ` �������P                           ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              �����������������������������������������������������                        �8   A �����@   ������   A �����@   �������@                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ����������?������������������������?�������������������                        8   �����@p   ������   �����@p   �������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ������������?�����������������������?����������������                        9�� ~?����[� � ��������� ~?����[� � ���������                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �7���?�����������������y�����?�����������������y����                        #9���~?����]�  ���������~?����]�  �������0                           ?�������     �������     �������     �������     �                           ��     �     �     8          �     �     8                             �{���������ƿ�����������k����������ƿ�����������k����                        9�� � ����X� P �������� � ����X� P �������                           ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8     D                        ����������?������������w���������?������������w����                        8 � �����@p >  ������ � �����@p >  �������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��7��������������������������������������������������                        �8 � ��?��@  |  W������ � ��?��@  |  W�������                            ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              �����������������������?�����������������������?���
��                         8����?��@ x������������?��@ x���������                            ?�������     �������     �������     �������     �                           @N     �     �     8          �     �     8                             �ݷ������}��������������������}����������������                        8��x���G����׀������x���G����׀�����                            ?�������     �������     �������     �������     �                           "N     �     �     8          �     �     8     $                        ��� ��������� >�����}��� ��������� >�����}����x                        A9���� @ �?��_���  � �������� @ �?��_���  � �����                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        ��6  ���������� ���������  ���������� �����������                        9����   0?��_���`  �������   0?��_���`  ����                           ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              ����  ����������  ����������  ����������  �����������                        )9����    ?��_���    �������    ?��_���    ����                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��7�  ����������  ����������  ����������  �����������                        9��� p  ?��W���    ������ p  ?��W���    ����                            ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              ����  ���������� ���������  ���������� ����������                        9���� 6  ?��_���` ` ������� 6  ?��_���` ` ����@                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      $                        �������������������������������������������������������                        8           @                     @          �@                           ?���������������������������������������������������                            O��������������������������������������������������                         ���                                                 ��                        b;���������������������������������������������������                            ?���������������������������������������������������                           O��������������������������������������������������                         ������������������������������������������������������                         8           @                     @          �                            ?���������������������������������������������������                           O��������������������������������������������������                        ������������c��!��/����;���������c��!��/����:��                        (9����� ?x�_�����`��������� ?x�_�����`�����                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                              ������������������]�/����8;���������������]�/����8:��                        9���>  ��_������ �������>  ��_������ �����                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��������������#���Yo�/����;�����������#���Yo�/����:��                         9��� � @��_������������ � @��_����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      D                        �6~� }r������`�/����:~� }r������`�/����:��                        .9������`A����_����8�����������`A����_����8�������                           >     �������     ?������     �������     ?�������                           ��     �     �     8          �     �     8                             ���>�,���x4������o���O�>�,���x4������o���O���                        ��������pA����_���>�����������pA����_���>������                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        ���>�r�,N���x4����/�������O�>�r�,N���x4����/�������O���                        �������p@����_���?<��������p@����_���?<���                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��7?��}#��߸�߳����>+����}�?��}#��߸�߳����>+����}���                         8��~��}p x��'O���-�� ��t��~��}p x��'O���-�� ��t�                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              �f�����r������?��(�����;����r������?��(�����:�h                         8/���o��E�B�������W��/���o��E�B�������W���                            >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     	�                        ������QB����믯���,���������QB����믯���,�������                        9�����  �P������  �������  �P������  ����                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8                             ��;�M�P�����������������
;�M�P�����������������
��                         ������ ���\�����
�������� ���\�����
����                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                             �߶38x�������3���?����38x�������3���?������                         9�����1����\�����W���������1����\�����W�����                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                             ��7���>���������������������>��������������������                        `8���?��@��@?����������?��@��@?��������                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              ������~ z�_�����/����u��������~ z�_�����/����u�������                        8��������A�������
���������A�������
��                            >     �������     ?������     �������     ?�������                           `N     �     �     8          �     �     8                             �������z�����������p���������z�����������p�������                         8?��w�}����A���������?��w�}����A����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      T                        ��63@�����/�����4���2�?���3@�����/�����4���2�?�����                         9̿�'�����\���������̿�'�����\����������                            >     �������     ?������     �������     ?�������                           @�     �     �     8          �     �     8                             ��a�����������{�?���a�����������{�?�����                         ����o�o����]� �����������o�o����]� ���������                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                             ���;��~������������ >��;��~������������ >����                        *9� ���q���_� ���������� ���q���_� ����������                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ������q�n�������XF����?�{���q�n�������XF����?�z��                        �9������ B����_������)��������� B����_������)����                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      D                        �����q������������o���?�;���q������������o���?�:�8                         9����� @��_�������������� @��_����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      �                        �߷���1�����������������?����1�����������������?���                        9����� @ ?��_�����P ������� @ ?��_�����P ���                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                             ��~����������������������
~����������������������
��                        9�����`@ ?�_���?� �������`@ ?�_���?� ����                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8                             �������������ƿ����h?����k����������ƿ����h?����j��                         8����~  �?@���?�� ������~  �?@���?�� ���                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��������������������?����J�����������������?����J�x                        �9�����~  �P������ �������~  �P������ ���`                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      �                        ������������������,��������������������,�������                         9�����~  ?�Q������� �������~  ?�Q������� ���                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ���o���������������������o�����������������������                        9������|  ?�Y������� � ������|  ?�Y������� � �                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                              ���������������������������������������������������                        9������8  � _�����Ӏ � ������8  � _�����Ӏ � �`                           >     �������     ?������     �������     ?�������                           PN     �     �     8          �     �     8                             �{���������������������������������������������������                         9������   � _������  � ������   � _������  � �                            >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     D                        ��7�����������������_������������������������_���������                        9������   @��_������  	�������   @��_������  	��                            >     �������     ?������     �������     ?�������                           `�     �     �     8          �     �     8                             ��������������������O������������������������O���������                         9������    ��_������   	�������    ��_������   	��                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              �����������������������������������������������������                        9������    �_������   �������    �_������   ��                            >     �������     ?������     �������     ?�������                           `N     �     �     8          �     �     8                             ��7�����~�����������������������~��������������������                         9������    ��_������   �������    ��_������   ��                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              �������~����������?������������~����������?����������                         9������   ? �_������  �������   ? �_������  ��                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              �������������������������������������������������������                        �������  � _������  � ������  � _������  � �                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                              �~7����������������������������������������������������                         9������   @ _������   ������   @ _������   �                            >     �������     ?������     �������     ?�������                           ��     �     �     8          �     �     8                             ������������������������������������������������������                        @9�������  @ _������   �������  @ _������   �                            >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8                             ��6G?�����?�����s���/������G?�����?�����s���/��������                        !9������o��@_������� < 5������o��@_������� < 4�                           >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              ���'?����?�����s�����������'?����?�����s������������x                        B9���?��w� x` _������ � ���?��w� x` _������ � �                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      �                        ���s����������;����������s����������;������������                        �������c� 9@ _������? � �����c� 9@ _������? � �                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        �����������������������������������������������������                        9������� �� _������ � ������� �� _������ � ��                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        ������?�����?������������������?�����?�����������������                        �9������ �� _������   ������ �� _������   �                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        ��������?������� /�����������?������� /��������                        �9��������_������� w���������_������� w��`                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��������������{�~/�����������������{�~/�������                        9�������^�������? `u�������^�������? `t�@                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8                             �n���}��� �?��������, ������}��� �?��������, ������                         9 ��������P >������ 5 ��������P >������ 4�                            >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     	                        �7��?y��� 0?��������� �����?y��� 0?��������� �����                        8  ������� @ ������   ������� @ ������ �                           >     �������     ?������     �������     ?�������                           ��     �     �     8          �     �     8                             ��������  ?���������  ��������  ?���������  �����                        �8�  ������  H  ������  �  ������  H  ������  �                            >     �������     ?������     �������     ?�������                           sN     �     �     8          �     �     8     4                        ��6������  ?���������  ���������  ?���������  �����                        9�  ���_���  \  ������  �  ���_���  \  ������  ��                           >     �������     ?������     �������     ?�������                           �     �     �     8          �     �     8     L                        ���'��i���  ?��������` ���'��i���  ?��������` �����                         ��  ������ M� ������X �  ������ M� ������X �                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                              ������������������������������������������������������x                        @8           @                     @          �                            ?���������������������������������������������������                           O�������������������������������������������������� �                        ���                                                 �x                         ;���������������������������������������������������                            ?���������������������������������������������������                           O�������������������������������������������������� �                        ������������������������������������������������������                         8           @                     @          �                            ?���������������������������������������������������                           �O��������������������������������������������������                        ���������������������������������������������                        $8 ���}����cA��������4 ���}����cA��������4�@                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �~7���>���w�|��������������>���w�|�������������                        @8  ��������@ �������84  ��������@ �������84�                            ?�������     �������     �������     �������     �                           ��     �     �     8          �     �     8                             ��7��� ����e����������[����� ����e����������[����                        8 ��}����#@��������4 ��}����#@��������4�                           ?�������     �������     �������     �������     �                           �     �     �     8          �     �     8                              �����������\�����8��������������\�����8�������                         9���������X��������5���������X��������4�                            ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8                             �������ꏾ������>���8|�[�����ꏾ������>���8|�Z��                        d9�������x4�\������O��������x4�\������O��@                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                             ���������������?(�����;������������?(�����:�h                        09������x4�\8��������O�������x4�\8��������O��                            ?�������     �������     �������     �������     �                           	N     �     �     8          �     �     8      �                        �_���~��~���_H�����-����u���~��~���_H�����-����u���                        D�����?�߸��\ 9�������}�����?�߸��\ 9�������}��H                           ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8     
                        ���/���o������������O���A�/���o������������O���A��h                         9��������_�`_�п����5��������_�`_�п����4�                            ?�������     �������     �������     �������     �                           	N     �     �     8          �     �     8      �                        ��7����������P����������E����������P����������E
��                        `9� ��A����_� ��������� ��A����_� ���������                            ?�������     �������     �������     �������     �                           �     �     �     8          �     �     8                             ���������S�?�����(��7�C��������S�?�����(��7�C���                        Q9����q�����_�+ ����������q�����_�+ �������                           ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8                             �۷��������~������h��y�G���������~������h��y�G���                         9�����s����_�~8��?���������s����_�~8��?�����                            ?�������     �������     �������     �������     �                           $N     �     �     8          �     �     8     D                        ������?���O��?����/���� z���?���O��?����/���� z��                        9���� �����_�<����������� �����_�<���������                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �۶������?_������������������?_��������������                        9�����_����_�p(�Pu����������_����_�p(�Pu������                           ?�������     �������     �������     �������     �                           $N     �     �     8          �     �     8     D                        ��?��w���@�������$�!�?��w���@�������$�!���                         9���������_o��Pp��������������_o��Pp������                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                             ���̿�'���<?�>���������c�̿�'���<?�>���������c���                        9����s/����_����W2�?�������s/����_����W2�?����                           ?�������     �������     �������     �������     �                           PN     �     �     8          �     �     8                             ������o��C�o�>�� ����?��C����o��C�o�>�� ����?��C���                        9���A�w����[����W{�?������A�w����[����W{�?����                            ?�������     �������     �������     �������     �                           @N     �     �     8          �     �     8                             �˷� ������_�f�� ��������Fk� ������_�f�� ��������Fj��                         ������e����\_���W� >�������e����\_���W� >���                           ?�������     �������     �������     �������     �                           4N     �     �     8          �     �     8     D                        ��7��������`y���������Ǒ���������`y���������Ǒ���                         8
�������@�������?�t
�������@�������?�t�                            ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              ���������������������9���������������������9�����                         8 q������@�����?�4 q������@�����?�4�                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      $                        �o7���������~>������o���������������~>������o��������                         8  �������@ �����?�  �������@ �����?��                            ?�������     �������     �������     �������     �                           ��     �     �     8          �     �     8     	                        �����������������?�)���w����������������?�)���w����                         9�  �������X ��������  �������X ��������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ����������������?����7���������������?����7����                        �9�  ~ ������_� ��?����e�  ~ ������_� ��?����d��                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                              �������ҽ���������+���������ҽ���������+�������                        9�  ~ }C�����_� ��?����E�  ~ }C�����_� ��?����D�@                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��7�������������������K�������������������J��                        9�  � mG�����_� ��������  � mG�����_� ���������                           ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              �����������������������������������������������x                        @9�  � g�����_  � V������  � g�����_  � V������                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        �������������������������������������������������                         8�  ~ �����N  � �������  ~ �����N  � �������                            ?�������     �������     �������     �������     �                           AN     �     �     8          �     �     8                             ���������������������������������������������������                         �   ~ �����@  � ������   ~ �����@  � �������                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��7����������a����������������������a��������������                         8  ~�����@  '�������  ~�����@  '��������                            ?�������     �������     �������     �������     �                           @�     �     �     8          �     �     8                             �������������a?����������������������a?��������������                         8   �����@   '�������   �����@   '��������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��������������?�����������������������?��������������                         �    �����@   �������    �����@   ��������                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                              ������������p����������������������p��������������                        C8   ?������@   #�������   ?������@   #��������0                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                             ���������������������������������������������������                        8   �������@  �8������   �������@  �8�������@                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      $                        ��7���������������������g�����������������������g���p                        �8@  f �����D  ` ������@  f �����D  ` �������                            ?�������     �������     �������     �������     �                           8�     �     �     8          �     �     8     �                        �����������������������������������������������������                        ��   A �����@   ������   A �����@   �������H                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ����������?������������������������?�������������������                         8   �����@p   ������   �����@p   �������                            ?�������     �������     �������     �������     �                           CN     �     �     8          �     �     8     4                        ������������?�����������������������?����������������                         9�� ~?����[� � ��������� ~?����[� � ��������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ������?�����������������y�����?�����������������y����                         9���~?����]�  ���������~?����]�  �������                            ?�������     �������     �������     �������     �                           AN     �     �     8          �     �     8                             ����������ƿ�����������k����������ƿ�����������k����                        9�� � ����X� P �������� � ����X� P �������                           ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8                             ����������?������������w���������?������������w����                         8 � �����@p >  ������ � �����@p >  �������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ����������������������������������������������������x                         8 � ��?��@  |  W������ � ��?��@  |  W�������                            ?�������     �������     �������     �������     �                           hN     �     �     8          �     �     8     �                        �����������������������?�����������������������?���
��                        8����?��@ x������������?��@ x���������                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ���������}��������������������}����������������                        8��x���G����׀������x���G����׀������                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ��� ��������� >�����}��� ��������� >�����}����x                        9���� @ �?��_���  � �������� @ �?��_���  � �����                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        ��  ���������� ���������  ���������� ����������8                         9����   0?��_���`  �������   0?��_���`  ����                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        ��6�  ����������  ����������  ����������  �����������                         9����    ?��_���    �������    ?��_���    ����                            ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              ��7�  ����������  ����������  ����������  �����������                         9��� p  ?��W���    ������ p  ?��W���    ����                            ?�������     �������     �������     �������     �                            �     �     �     8          �     �     8                              ����  ���������� ���������  ���������� ����������                         9���� 6  ?��_���` ` ������� 6  ?��_���` ` ����                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      $                        ��7���������������������������������������������������p                        �8           @                     @          �                            ?���������������������������������������������������                           ��������������������������������������������������� �                        ���                                                 ��                        ����������������������������������������������������                           ?���������������������������������������������������                            O��������������������������������������������������                         �Ϸ����������������������������������������������������                        ��           @                     @          �                           ?���������������������������������������������������                           0O��������������������������������������������������                        ��7���������c��!��/����;���������c��!��/����:��                        49����� ?x�_�����`��������� ?x�_�����`�����@                           >     �������     ?������     �������     ?�������                           �     �     �     8          �     �     8                              �޷���������������]�/����8;���������������]�/����8:��                        �����>  ��_������ �������>  ��_������ �����                           >     �������     ?������     �������     ?�������                           !N     �     �     8          �     �     8                             ��������������#���Yo�/����;�����������#���Yo�/����:�x                         9��� � @��_������������ � @��_����������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      �                        ��6~� }r������`�/����:~� }r������`�/����:��                         9������`A����_����8�����������`A����_����8������                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              ���>�,���x4������o���O�>�,���x4������o���O���                         9������pA����_���>�����������pA����_���>������                            >     �������     ?������     �������     ?�������                           PN     �     �     8          �     �     8                             ���>�r�,N���x4����/�������O�>�r�,N���x4����/�������O���                        P9������p@����_���?<��������p@����_���?<���                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��7?��}#��߸�߳����>+����}�?��}#��߸�߳����>+����}���                         8��~��}p x��'O���-�� ��t��~��}p x��'O���-�� ��t�                            >     �������     ?������     �������     ?�������                           P�     �     �     8          �     �     8                             �������r������?��(�����;����r������?��(�����:��                        �/���o��E�B�������W��/���o��E�B�������W���                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              �������QB����믯���,���������QB����믯���,�������                         9�����  �P������  �������  �P������  ���                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ���;�M�P�����������������
;�M�P�����������������
��                        9����� ���\�����
�������� ���\�����
����                           >     �������     ?������     �������     ?�������                           @N     �     �     8          �     �     8                             ���38x�������3���?����38x�������3���?������                        �9�����1����\�����W���������1����\�����W�����                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ������>���������������������>��������������������                         8���?��@��@?����������?��@��@?��������                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      D                        ������~ z�_�����/����u��������~ z�_�����/����u�������                        @8��������A�������
���������A�������
��                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              �?7����z�����������p���������z�����������p�������                        8?��w�}����A���������?��w�}����A����������                           >     �������     ?������     �������     ?�������                           ��     �     �     8          �     �     8                             ��63@�����/�����4���2�?���3@�����/�����4���2�?�����                        �9̿�'�����\���������̿�'�����\����������                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              ���a�����������{�?���a�����������{�?�����                        9���o�o����]� �����������o�o����]� ���������                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              �۶;��~������������ >��;��~������������ >����                        9� ���q���_� ���������� ���q���_� ����������                            >     �������     ?������     �������     ?�������                           $N     �     �     8          �     �     8     D                        ������q�n�������XF����?�{���q�n�������XF����?�z��                         9������ B����_������)��������� B����_������)����                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      D                        ��7���q������������o���?�;���q������������o���?�:��                        9����� @��_�������������� @��_����������@                           >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              ��7���1�����������������?����1�����������������?��`                        9����� @ ?��_�����P ������� @ ?��_�����P ���                            >     �������     ?������     �������     ?�������                           	�     �     �     8          �     �     8      �                        ��6~����������������������
~����������������������
��                        9�����`@ ?�_���?� �������`@ ?�_���?� ���@                           >     �������     ?������     �������     ?�������                           A�     �     �     8          �     �     8                             �������������ƿ����h?����k����������ƿ����h?����j��                        8����~  �?@���?�� ������~  �?@���?�� ���                           >     �������     ?������     �������     ?�������                           bN     �     �     8          �     �     8     $                        ��6�����������������?����J�����������������?����J��                         9�����~  �P������ �������~  �P������ ���                            >     �������     ?������     �������     ?�������                           �     �     �     8          �     �     8      ,                        ������������������,��������������������,�������                         9�����~  ?�Q������� �������~  ?�Q������� ���                            >     �������     ?������     �������     ?�������                           dN     �     �     8          �     �     8     D                        ���o���������������������o�����������������������                         9������|  ?�Y������� � ������|  ?�Y������� � �                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        ���������������������������������������������������                        �9������8  � _�����Ӏ � ������8  � _�����Ӏ � �                            >     �������     ?������     �������     ?�������                           QN     �     �     8          �     �     8                             �����������������������������������������������������                        �9������   � _������  � ������   � _������  � ��                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��������������������_������������������������_��������x                        �9������   @��_������  	�������   @��_������  	��                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      �                        �������������������O������������������������O���������                        9������    ��_������   	�������    ��_������   	��`                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8                             �����������������������������������������������������                        9������    �_������   �������    �_������   ��                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��������~�����������������������~��������������������                        �9������    ��_������   �������    ��_������   ��                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        �������~����������?������������~����������?����������                        9������   ? �_������  �������   ? �_������  ��@                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      $                        �������������������������������������������������������                         �������  � _������  � ������  � _������  � �                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8      T                        �������������������������������������������������������                        �������   @ _������   ������   @ _������   �(                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��7����������������������������������������������������                        "9�������  @ _������   �������  @ _������   �                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                              ��6G?�����?�����s���/������G?�����?�����s���/��������                         9������o��@_������� < 5������o��@_������� < 4�                            >     �������     ?������     �������     ?�������                           �     �     �     8          �     �     8      ,                        ���'?����?�����s�����������'?����?�����s�������������                         9���?��w� x` _������ � ���?��w� x` _������ � �                            >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ��6s����������;����������s����������;������������                        �9�����c� 9@ _������? � �����c� 9@ _������? � �                            >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                             �����������������������������������������������������                        f9������� �� _������ � ������� �� _������ � �`                           >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          