�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������_���������������������������������_���������������������������������_�������������������������������?�����������������������������������_���������������������������������_���������������������������������_�������������������������������?�����������������������������������Og�0�&4�1��>�����Ɵm������������Og�0�&4�1��>�����Ɵm������������Og�0�&4�1��>�����Ɵm����������?�����������������������������������_[��]o�_n��uޛ�S]�omu������������_[��]o�_n��uޛ�S]�omu������������_[��]o�_n��uޛ�S]�omu����������?�����������������������������������_o��]n_n��޻�W]ꮂ�Uu������������_o��]n_n��޻�W]ꮂ�Uu������������_o��]n_n��޻�W]ꮂ�Uu����������?�����������������������������������_w��]m�_n��}޻�W]ꮾ�Uu������������_w��]m�_n��}޻�W]ꮾ�Uu������������_w��]m�_n��}޻�W]ꮾ�Uu����������?�����������������������������������_[��]m�_n��u޻�W]�n��u������������_[��]m�_n��u޻�W]�n��u������������_[��]m�_n��u޻�W]�n��u����������?�����������������������������������og���vo��c�>��Wa�n�ﻍ�����������og���vo��c�>��Wa�n�ﻍ�����������og���vo��c�>��Wa�n�ﻍ���������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������o�������������������������������o�������������������������������o�����������������������������?�����������������������������������o�������������������������������o�������������������������������o�����������������������������?�����������������������������������)�}���1��.ƶ�Lm�p�~bq�&18���������)�}���1��.ƶ�Lm�p�~bq�&18���������)�}���1��.ƶ�Lm�p�~bq�&18�������?�����������������������������������f�����n�]n���_����k����o����������f�����n�]n���_����k����o����������f�����n�]n���_����k����o��������?�����������������������������������n�����`�_n¶�\*����>�n���������n�����`�_n¶�\*����>�n���������n�����`�_n¶�\*����>�n�������?�����������������������������������n�����o�_n���[������m��m�����������n�����o�_n���[������m��m�����������n�����o�_n���[������m��m���������?�����������������������������������n��n��n�]l���[�k��뽭��m����������n��n��n�]l���[�k��뽭��m����������n��n��n�]l���[�k��뽭��m��������?�������������������������������������~���q�c�»�\7k���~m��n������������~���q�c�»�\7k���~m��n������������~���q�c�»�\7k���~m��n��������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������>S����q�S���c�p���N>�o�����������>S����q�S���c�p���N>�o�����������>S����q�S���c�p���N>�o��������?�����������������������������������t��w������w��]�o���{5���_����������t��w������w��]�o���{5���_����������t��w������w��]�o���{5���_��������?�����������������������������������u����������A�l.��{t��?����������u����������A�l.��{t��?����������u����������A�l.��{t��?��������?�����������������������������������u����������_�k���{u���_����������u����������_�k���{u���_����������u����������_�k���{u���_��������?�����������������������������������u��w������w��]�k���{u�v�o����������u��w������w��]�k���{u�v�o����������u��w������w��]�k���{u�v�o��������?�������������������������������������]���{��]���c�l0��}v?ww������������]���{��]���c�l0��}v?ww������������]���{��]���c�l0��}v?ww��������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?��������������������������������������Ɍ��&5?q��s��c0��1�������������Ɍ��&5?q��s��c0��1�������������Ɍ��&5?q��s��c0��1��������?����������������������������������������u�]o��뮿Z����}n��~���������������u�]o��뮿Z����}n��~���������������u�]o��뮿Z����}n��~��������?�����������������������������������������n�렸Z���an��p����������������n�렸Z���an��p����������������n�렸Z���an��p��������?�����������������������������������u����}��m��믷Z����]n��n����������u����}��m��믷Z����]n��n����������u����}��m��믷Z����]n��n��������?�����������������������������������u���[u�]m��뮷Z����]n��nݮ��������u���[u�]m��뮷Z����]n��nݮ��������u���[u�]m��뮷Z����]n��nݮ������?��������������������������������������]���v�q�k���ap��pݮ�����������]���v�q�k���ap��pݮ�����������]���v�q�k���ap��pݮ������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������W����������������������������������W����������������������������������W����������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������mW͵1�ɌO��lev6�f5������������mW͵1�ɌO��lev6�f5������������mW͵1�ɌO��lev6�f5��������?��������������������������������������mW��n��u��ۯ�u����u޶������������mW��n��u��ۯ�u����u޶������������mW��n��u��ۯ�u����u޶�������?�������������������������������������UW�Uo��u���,-���.޶��?���������UW�Uo��u���,-���.޶��?���������UW�Uo��u���,-���.޶��?�����?�����������������������������������u��UW�Uo��u���뭭�����}޶����������u��UW�Uo��u���뭭�����}޶����������u��UW�Uo��u���뭭�����}޶��������?�����������������������������������u��W��n��u��۫���>��u޶���������u��W��n��u��۫���>��u޶���������u��W��n��u��۫���>��u޶�������?��������������������������������������W��ۍ���l5�7v�������������W��ۍ���l5�7v�������������W��ۍ���l5�7v��������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������{���������������������������������{���������������������������������{�����������������������?�����������������������������������������������o��������������������������������o��������������������������������o������������������?�����������������������������������������������o�������������������������������o�������������������������������o�����������������?�����������������������������������1���p��8z'1��)�ɌN?�sS�����������1���p��8z'1��)�ɌN?�sS�����������1���p��8z'1��)�ɌN?�sS���������?�����������������������������������n�{o����z���_f�����ݯ�Mw����������n�{o����z���_f�����ݯ�Mw����������n�{o����z���_f�����ݯ�Mw��������?�����������������������������������n�{l.��z���_n�ۅ�ݬ7]w����������n�{l.��z���_n�ۅ�ݬ7]w����������n�{l.��z���_n�ۅ�ݬ7]w��������?�����������������������������������n�{k����z���_n��u�����]w����������n�{k����z���_n��u�����]w����������n�{k����z���_n��u�����]w��������?�����������������������������������n�{k����z���_n��u�߾��]wݫ��������n�{k����z���_n��u�߾��]wݫ��������n�{k����z���_n��u�߾��]wݫ������?�������������������������������������{l0��8z�1�߮�ۅ�7��3]�ݫ����������{l0��8z�1�߮�ۅ�7��3]�ݫ����������{l0��8z�1�߮�ۅ�7��3]�ݫ������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������������������߂��������������������������������߂��������������������������������߂����������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������8����c�Ӎ���>ϧ������������8����c�Ӎ���>ϧ������������8����c�Ӎ���>ϧ����������?�����������������������������������u�]mw����Mu�]u��j޷��m������������u�]mw����Mu�]u��j޷��m������������u�]mw����Mu�]u��j޷��m����������?�����������������������������������t�m����]u�_���~ߺ�m������������t�m����]u�_���~ߺ�m������������t�m����]u�_���~ߺ�m����������?�����������������������������������u��m����]u�_}�����mu�����������u��m����]u�_}�����mu�����������u��m����]u�_}�����mu���������?�����������������������������������u�]mw����]u�]u���޷��mu�����������u�]mw����]u�]u���޷��mu�����������u�]mw����]u�]u���޷��mu���������?�����������������������������������8�m�����ݎWc���>ϻm�����������8�m�����ݎWc���>ϻm�����������8�m�����ݎWc���>ϻm���������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        