�P��<o ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                               ��                               ��                               ��                               ��                               ��                               ��                               ��              ����������������@��0  ? `                       ���0  ? `                       ���0  ? `                       ���0  ? `                       @��0 1�`�                     s���0 1�`�                     s���0 1�`�                     s���0 1�`�    ����������������@� 0 1�`�                     y�� 0 1�`�                     y�� 0 1�`�                     y�� 0 1�`�                     @�3ǜ1�g��                     |��3ǜ1�g��                     |��3ǜ1�g��                     |��3ǜ1�g��    ����������������@���l�?lٙ�                    ~>���l�?lٙ�                    ~>���l�?lٙ�                    ~>���l�?lٙ�                    @� ߷�0oٟ�                    ~>� ߷�0oٟ�                    ~>� ߷�0oٟ�                    ~>� ߷�0oٟ�   ����������������@� �603l�                     |�� �603l�                     |�� �603l�                     |�� �603l�                     @�ٶl�03lٙ�                    y��ٶl�03lٙ�                    y��ٶl�03lٙ�                    y��ٶl�03lٙ�   ����������������@��3ǌ0g��                     s���3ǌ0g��                     s���3ǌ0g��                     s���3ǌ0g��                     @�                               ��                               ��                               ��              ����������������@�                               ��                               ��                               ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����xq�������������������������������xq�������������������������������xq����������������������������                                 ���������_�������������������������������_�������������������������������_�����������������������                                 ����ׯ����_���������������������������ׯ����_���������������������������ׯ����_������������������������ >          �         �         ����ׯ����O�����v�8��������cg����������ׯ����O�����v�8��������cg����������ׯ����O�����v�8��������cg������� "          �                   ����ױ���]_����_���W�������[����������ױ���]_����_���W�������[����������ױ���]_����_���W�������[������� "          �                   ����׾���]_����\6��P�������o����������׾���]_����\6��P�������o����������׾���]_����\6��P�������o������� "          �                   ����׾���]_����[���W��������w����������׾���]_����[���W��������w����������׾���]_����[���W��������w������� >          �         �         �������n�Y_����[���W�������[�������������n�Y_����[���W�������[�������������n�Y_����[���W�������[�������                                 ����xq��eo����\;�8X�������ag����������xq��eo����\;�8X�������ag����������xq��eo����\;�8X�������ag�������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����?����������o����������������������?����������o����������������������?����������o�������������������                                 ���������������_{�����������_��������������������_{�����������_��������������������_{�����������_������                                 ���������������_�����������_��������������������_�����������_��������������������_�����������_������ >          �         �         �������?������cO~c��������8Ͽ������������?������cO~c��������8Ͽ������������?������cO~c��������8Ͽ������ "          �                   �������������}_b����������_�������������������}_b����������_�������������������}_b����������_������� "          �                   �������������aYz���������_W������������������aYz���������_W������������������aYz���������_W������ "          �                   �������������]_zݷ������u��o������������������]_zݷ������u��o������������������]_zݷ������u��o������ >          �         �         ������n��������]_r��������u�_o�����������n��������]_r��������u�_o�����������n��������]_r��������u�_o������                                 ����7�?������a_����������8ߗ���������7�?������a_����������8ߗ���������7�?������a_����������8ߗ������                                 ����������������������������������������������������������������������������������������������������������                                 �������������������?����������������������������������?����������������������������������?����������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����?���������o���������������������?���������o���������������������?���������o������������������                                 ��������������_u�������������������������������_u�������������������������������_u������������������                                 ��������������_u�������������������������������_u�������������������������������_u������������������ >          �         �         ������cg�������cOuv?�������q�������������cg�������cOuv?�������q�������������cg�������cOuv?�������q�������� "          �                   ����?Z�[�������}_u�������ۮ�����������?Z�[�������}_u�������ۮ�����������?Z�[�������}_u�������ۮ�������� "          �                   �����n�o�������aYut�����껮������������n�o�������aYut�����껮������������n�o�������aYut�����껮�������� "          �                   �����v�w�������]_uu������껮������������v�w�������]_uu������껮������������v�w�������]_uu������껮�������� >          �         �         �����Z�[�������]_ue�������{�������������Z�[�������]_ue�������{�������������Z�[�������]_ue�������{���������                                 �����gcg�������a_�?������|q������������gcg�������a_�?������|q������������gcg�������a_�?������|q��������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����/����������o}�������������������/����������o}�������������������/����������o}����������������                                 ���������������_}������������������������������_}������������������������������_}����������������                                 ���������������_�������������������������������_�������������������������������_����������������� >          �         �         �����f7��������cO�cc?������0������������f7��������cO�cc?������0������������f7��������cO�cc?������0�������� "          �                   ����k����������}_�]]�����u�W���������k����������}_�]]�����u�W���������k����������}_�]]�����u�W������ "          �                   �������������aY�]A������P������������������aY�]A������P������������������aY�]A������P������ "          �                   ��������������]_�]_�����}�W��������������������]_�]_�����}�W��������������������]_�]_�����}�W������� >          �         �         ��������������]_�]]�����u�W�������������������]_�]]�����u�W�������������������]_�]]�����u�W������                                 �����n��������a_�cc�������0������������n��������a_�cc�������0������������n��������a_�cc�������0��������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ���������������o��������������������������������o��������������������������������o������������������                                 ���������������_w��������������������������������_w��������������������������������_w������������������                                 ���������������_w��������������������������������_w��������������������������������_w������������������ >          �         �         �����˦?�������cOv6�������c6�����������˦?�������cOv6�������c6�����������˦?�������cOv6�������c6������� "          �                   �����[���������}_���������v�����������[���������}_���������v�����������[���������}_���������v������� "          �                   ����X[��������aYt��������v����������X[��������aYt��������v����������X[��������aYt��������v������� "          �                   �����[���������]_u����������v�����������[���������]_u����������v�����������[���������]_u����������v������� >          �         �         �����[-��������]_u���������y�����������[-��������]_u���������y�����������[-��������]_u���������y�������                                 �����l�?�������a_6�������a{�����������l�?�������a_6�������a{�����������l�?�������a_6�������a{�������                                 ����������������������������������������������������������������������������������������������������������                                 �������������������?����������������������������������?����������������������������������?����������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������