�P   ˀ�                                                                                                                                                                 ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                       ��                      �������������������������������������������������������� ?������������������������������������������������������������������������������������������������������                                                                                                                                       ��                      �������������������������������������������������������� ?������������������������������������������������������������������������������������������������������                                                                                                                                       ��                      �������������������������������������������������������� ?������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������                          ������������               ��        �����          ���������������������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������                          ������������               ��        �����          ���������������������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������         �                ������������               ��        �����          ���������?�����������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������         �                ������������               ��        �����          ���������?�����������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������         �                ������������               ��        �����          ���������?�����������������           �����������������������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ������������������������������� ������������������                         ��                                ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ������������������������������� ������������������                         ��                                ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ������������������������������� ������������������                         ��                                ��                 ?����������������������������������������������������������� ������������������                                                                                �������������������������� ����������������������������������������������������                         ��                                                   ?��������������������������������������������������������������������������������                                                                                �������������������������� ����������������������������������������������������                         ��                                                   ?��������������������������������������������������������������������������������                                                                                �������������������������� ����������������������������������������������������                         ��                                                    ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                               ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������          ��                                                                    �������������������������������������������������������������������������������                                                                                ���������� �������������������������������������������������������������������          ��                                                                    �������������������������������������������������������������������������������                                                                                ���������� �������������������������������������������������������������������   �      ��                                                                   ������������������������������������������������������ �����������������������   �                                                                           ��������� ������������������������������������������ �����������������������  �      ��                                                                   ������������������������������������������������������ �����������������������  �                                                                           ���?������ ������������������������������������������ �����������������������  �      ��                                                                �  ������������������������������������������������������ ����������������������  �                                                                        �  ���_������ ������������������������������������������ ��������������������?��  �      ��                                                                �  ����?������������������������������������������������� ����������������������  �                                                                        �  ���?������ ������������������������������������������ ����������������������  ?�      ��                                                                �  ����������������������������������������������������� ����������������������  ?�                                                                        �  ��������� ������������������������������������������ ����������������������  x      ��                                                               �<  ����������������������������������������������������� ����������������������  x                                                                          <  ��������� ������������������������������������������ ����������������������  ��      ��               �������������������������                       �  ����������������������������������������������������� ����������������������  ��                       �������������������������                       �  �������� ������������������������������������������ ��������������������!�� �@     ��               ?�������������������������                      �_  ��������� ������������������������������������������ ����������������������� �      ��               ?�������������������������                      �K  �������� ���������������                        �� �������������������� �� �@     ��               �������������������������                      �  �������� ������������������������������������������ �����������������������        ��               �������������������������                      �  ��(������ ���������������                        �� ��������������������(�� ��      ��               ��������������������������                       Ӏ ��������� ���������������?�������������������������� ������������������ ��� ��      ��               �?������������������������                       Ӏ ��h������ ����������������                      �� ��������������������,� �      ��              ��������������������������                      �� ���]����� ����������������������������������������� ������������������t?���         ��              �������������������������~                         � ��(������ ��������������                        ��� ��������������������(� �  @                    ��                      �                       � ��'�^�������������������������������������������������� ���������������������o�                          ��������������������������                        @ �� �����������������������                      @A�� ������������������
  ?� ��                      ��         ���         ��                       �� ��?� ?�����������������������                     ��� ������������������ ��� ?�                       ��                     �                       �� �������������������������� �����������������������!�� ��������������������� �                       ��������������������������                        ?� ��/�^������������������������������������������������������������������������� (                        �������������������������                        (P ��  �����������������������          @            �!����������������������
  /� �                       �������������������������                        � ��+�^�������������������������������������������������������������������������� (                        ��������������������������                        (P ��  �����������������������           @             ����������������������
  /� ��                      �������������������������                       �� ��� ?��������������������������������������������������������������������� ��� �                       ��������������������������                       �� ��������������������������           @             ������������������������� �                      ��         8           �                      � �� ��)�\����������������������������������������������������������������������u�(� (                        ������������  �����������                        (@ ��  �����������������������           @             ����������������������
  ?� �                      ��         ;���         ?�                      ��� ��(�X������������������������         <  >         �����������������������5�(� (                        ��         8           �                        (@ ��  ����������������������� ����������  !��������������������������������
  ?� ��\                     �������������������������|                      t�� ��(? ���������������������������������  ?����������������������������������(�� ~(                        ������������  �����������                        (� ��  �����������������������           @             �����������������������  � �                     �?������������������������                     ���� ������������������������������������  ?�������������������������������������� �                      ������������  �����������                     ���� ��� �����������������������           @             ����������������������> � ��         ��������������������������������������������������          ?�0 ����?���������            ������������  ?�����������           �����������?� ��                      ������������  �����������                     �0 �������������������������           @             �������������������������� ���         �������������          ;���          ?������������          ?��p ��(��?���������������������������������  ?����������������������������������*)�� (��         ������������������������ 0�����������������������          
*)p ��  ����������                       @ 0                        �����������  �� ���         �������������          ;���          ?������������          ��0 �����?����������������������          < 0>          ?�����������������������+�� ���         �������������          8 p          ?�������������         
*0 �� (����������            ����������� 0!�����������            ����������(���������       ���������������������������������������������������       ������      �������������������������������� p?�������������������������������                   ������������������������ p�����������������������             ���������������|                      @ p                      �?���������������������       ��������������������������������������������������       ?���������������������}����������������������� �?���������������������������������������������       }����������������������� �������������������������       ?������      ���������                      @ �                      ��������      �������       ��������������������������������������������������       ����������������������������������������������?���������������������������������������������       �������������������������������������������������       ������      ��������                      @�                      ��������      �������       ��                     ;�/�                     ��       ����������������������������������������������?���������������������������������������������       ������������������������������������������������       �������       �������� �                     @�                      ��������      �������       ��                     ;�O�                     ��      �����������������������                      <�>                     ������������������������      �                      8�                     ��       �������       ������� ������������������������!�����������������������������       �������       �������������������������������������������������      ����������������������������������������������`?����������������������������������������������      ������������������������;�������������������������       �������       �������                       @?`                        �������       �������       ������������������������?�������������������������      �����������������������������������������������?����������������������������������������������      ������������������������ ������������������������       �������       �������                       @�                        �������       �������       ����������������  ����������  ?�����������������      ����������������������������������������������?�?����������������������������������������������      ������������������������  ������������������������       �������       �������                       @?�                        �������       �            ����������������     ;���   0  �����������������      �     ��������������������������������������� ?����������������������������������������������      �����������������  ����  ����  ?�����������������       �������       �������                 ���   @     ���                �������       �            |���������������     ;���   0  �����������������      �     ��������������������������������   <  >   ?��������������������������������������      ����������������     8     8  ?�����������������       ������   ���������               �������  !�������              |��������   ���   ?�       �����������������  �����������  ����������������      ��   ���   ���������������������������������  ?���������������������������������   ���   ��      �����������������  ����  ����  ?�����������������       ��   �       �������                 ���   @      ���                �������      ��   ?����������������{����{����  ����  ����  ����{����{����������������   ���   ��      �������{����{�������������������������{����{�������      ��   ���   ��      �������{����{����  ����  ����  ?����{����{�������      ��   �       �������   !B�!B�!B ���   G���   ��� B�!B�!B   �������      ��   ?����������������{����{���������������8�����{����{����������������   ���   ����������������{����{������������������������{����{����������������   ���   ����������������{����{���������������8�?����{����{����������������   �                  !B�!B�!B ���   @      ��� B�!B�!B                 �     �������� �����{����{�����   ?���   0E����{����{��������������    ��   ����������������{����{�����]������������������{����{����������������   ���   ����������������{����{����������������E?����{����{����������������   �                  !B�!B�!B ���   @      ��� B�!B�!B                 �     �������� �����{����{�����   ?���   0E����{����{��������������    �    �������� �����{����{�����]�   ?���   ?������{����{��������������    �    �������� �����{����{�����   ?���   8E?����{����{��������������    �   ?�        �� !B�!B�!B �������  ������� B�!B�!B �        �   ���   ?��������������������������������������E��������������������������   ���   ���������������������������]����������������������������������������   ���   ��������������������������������������E?��������������������������   �                                ���   @      ���                              ��   ?������������             �����  ����E�            ������������   ���   ���������������������������]����������������������������������������   ���   �������������������������������  ����E?��������������������������   �                                ���   ���   ���                �             �� 0 ?������������             ������������E�            ������������  ���   ���������������������������]����������������������������������������   ��� 0 ������������             ������������E?�            ������������  �   0    ��    �����������������          ���������������� ����  p    �      ww�0?  ����������������          0E�����������������w|�  ?���   ������������             �]���������������            ������������   ���  ������������             ������������E?�            ������������ ?��       ww�0?   �����������������          ���������������� ��w|�  ?� �  �    |7�p  ����������������          0E������������������~�  ��      }��p  ����������������]�          ?����������������������    � �    |7�p  ����������������          8E?������������������~� � � � ?�����������               �����������������              ����������� ����� ?�������������������������������������8��������������������������� �����   ��������������������������������������������������������������������   ���� �������������������������������������8�?�������������������������� ���  �   ����                  ���          ���               ��w�~�  �� ��À?����������������{����{����  �����������  ����{����{�������?�����o� �����   ����������������{����{�������������������������{����{����������������   ���À����������������{����{����  �����������  ?����{����{�������?�����o� ���  À  �?���    !B�!B�!B ���          ��� B�!B�!B  �����  �� ��� ?������ϑ��������{����{����  �����������  ����{����{��������]����������   ����������������{����{�������������������������{����{����������������   ���� ������ϑ��������{����{����  �����������  ?����{����{��������]��������  �   >9�9���    !B�!B�!B ���          ��� B�!B�!B  ���?�>� �� � �   <y�1��� �����{����{����            0  ����{����{������<>�p À��   ����������������{����{�������������������������{����{����������������   ���� �������9��������{����{����  �����������  ?����{����{���������?�����À�  �   >y�9����   !B�!B�!B ���          ��� B�!B�!B  ��>�|| À �    <��a��� �����{����{����            0  ����{����{�����;<8>��< ���     <��q�σ� �����{����{�������          ?�������{����{�����?�<>��<    �   <��a��� �����{����{����            8  ?����{����{�����;<8>��<�� � ?����������� !B�!B�!B ����������������� B�!B�!B ���������������� ?��?� p�?���������������������������������������������������C�À �������   ��<?�`q������������������  �����������  ?������������������ǀ��   ��� ��?� p�?�����������������  �����������  ?�����������������C�À �����     }��w���                 ���          ���               �<���< �� �� ?��? p�?����������������������������������������������������ǀ��������   ��<@q�����������������������      �����������������������ǀ���   ��� ��? p�?����������������������      �����������������������ǀ������     ������                     ?�������                    <8?��| �� �� ?��>@q��������������������������������������������������� ��� �� ���   ��~|�������������������������������������������������������� ��   ��� ��>@q��������������������������������������������������� ��� �� �     ��翎�                                                 �<8����� �  �� ?��8<@q���������������������������������������������������Ã� ��� ���   ��8�������������������������������������������������������yÏ���   ��� ��8<@q���������������������������������������������������Ã� ��� �     ��ÿ�?�        |                                �      �<|9�;��� �  ��< ?��|�����������������������������������������������������'� ��� ���   ����������������������������������������������������������?�qϏ��   ���< ��|�����������������������������������������������������'� ��� �  <   ���?�        @                                �      �?�;�3��� �  ��� ?����� ������������������������������������������������������� �� ���   ��������������������������������������������������������������ρ��   ���� ����� ������������������������������������������������������� �� �  �   ~���         @             !<�x           � �      �?p?�q��� �  ��   ?�� ��������������������������������������������������������?�q����   ���   �������������������������������������������������������������������   ���   �� ��������������������������������������������������������?�q����   �       |��w         @�q�          1B�D           ��       ~?�;�pp�p     ��   ?��������������������������������������������������������������ρ��   ���   ���������������������������������������������������������������������   ���   ��������������������������������������������������������������ρ��   �       8��         y�           1BD�B           L��       | p0~p     ��   ?�������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   �������������������������������������������������������������������   �                   A��          )BD�B           H��       0   `` `     ��   ?���������������������������������������������������������������������   ���   �������������������}�����������������������������7]_�����������������   ���   �������������������}�����������������������������7]_�����������������   �                      A�           )BD�B           Ȣ�               `     ��   ?���   �������������������������������������������������������   ����   ���   �������������������u�����������ڽ�WZ��������������]]�����������������   ���   �������������������u�����������ڽ�WZ��������������]]�����������������   �                       A�           %B��B           (��                     ��   ?���������������������������������������������������������������������   ���   �������������������?����������ܽ�W\��������������ac�����������������   ���   �������������������?����������ܽ�W\��������������ac�����������������   �                      @�q�          #B��B           (��                    ��   ?���   �������������������������������������������������������  ����   ���   �������������������������������ܽ��\���������������������������������   ���   ���   ������������������������ܽ��\��������������������������  ����   �         ����                        #B�D                       ���        ��   ?��������������������������������������������������������������������   ���   �����������������������������������^���������������������������������   ���   ����������������������������������^���������������������������������   �         �  (                        !<�x             <                    ���������������������������������������������������������������������������������   ���������������������������������������������������������������������   ���   ��������������������������������������������������������������������   � ����   �  (                                                           ���� ���������   �������������������������������������������������������  ������������������   �������������������������������������������������������  ������������������   �������������������������������������������������������  ���������         ����                                                      ���         ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ���������   ������������������������      ������������������������   ������������������   �������������������������������������������������������   ������������������   �������������������������������������������������������   ���������        ����                                                      ?���         �������������������������������������      ���������������������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������������                                    ?�������                                    ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            