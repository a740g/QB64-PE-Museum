�P   ˀ� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                <x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �` �0 �  `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                          ` �                                                                           ` �                                    0 �   `   `� � 8 ό 8 ` � p�p��q�� |��9� �   0 �   `   ���������������������������������������������������������?����������������                  `` �  �  8    � p`p��p3� ��9�                                     `` �  �  8    � p`p��p3� ��9�                      0 �   `   ��� ����� ` ���s������� ||ws�w�0?�   0 �   `   ������������������������������������������������������������?����������������                 ��� �����    ��xs������� |<wp�w�0?                                   ��� �����    ��xs������� |<wp�w�0?                     0 �   `   �?�� ���� ` ���v<����`< 8x|3�w�p�   0 �   `   �������������������������������������������������������������?����������������                 �?�� ����    ���v<����`< 88|1�w�p                                   �?�� ����    ���v>À��`< <8|1�w�p                     0 �   `   �<�<?� �ǁ��p ` ���p8�� ��px �x�;������   0 �   `   ������������������������������������������������������������?����������������                 �<8<;� �ǁ��p    ���p8�� ��px �8�;�����                                   �>x<;� �����x    ���p>�����~ �<�������                    0 �   `   �<<8q� ��Ǉ0 ` �c�x8� ��p� ���?������   0 �  a_  ������������������������������������������������������������?����������������               �<<8q� ��Ǉ0    �c8x8� ��p� ���?�����            A_                  �?�<� �ϻ����    ��x{�������� ��������            A_     p �   `   �|~p� ����  � ��8 8�r���a� p��3���À�   0 �  aD  �������������������������������������������������������������?����������������   @           �|~p� ����  � ��8 8�p���a� p��1���À            AD      @           ��|�����ϟ� � ��?���|����a� x��1�����            AD     p �   `   ����p����8 ���p9�v�c��c�����3�����   0 �  bD  �����������������������������������������������������������������������������   @           �~��p����8 ���p9�p�c��c�����3�����           "D      @           �<~����ρ�߿~ ����~���x��c��s�����;������           "D    
�}���  `   �8�c����x��?��<���;0a��Ï ��c�����   0 �  tD  ����������������������������������������������������������������������������  
�m�r�        �8c����x��?��<w��; a��Ï ��c�����           D     
�m�r�        �<{������~>��?�����?�a���� ���������           D    )yS�)  `                       �   0              @   0 �  hD  ������������������G�y �������|�`��?�ώx8���?�x `q�?����������������  )IR�)                                                                 D     )IR�)        �}���������|�����8|���q���� ���s���σ�           D    
$y�$  `                       �   0                  0 �  tD  ��������������������x� ������`��@��>�����p�<x@q�����������������  
$I�$                                                                 D     
$I�$        �8��������x>����|y��o�s�������������           D      0     `             �              0                   0 �   @   ���݆��u������������0<x� ��f������<9������x ~|p����������������                                                                                  
"I�"        �x������x����<������ ��Ϗ���������           "D      0     `             �              0               @   0 �       ���ֆˬu����������!�8<p?�a�g���|�!<8xy���q�����8�`�����������������                                                                                  
)I4R�)        �=������;<�q����������� ���~ �s�c����?�           AD       �   `           �               0               @   0 �       �����,t����������a�><a?�`gǀg��<�0c�<>����������G������������������                                                                                  
&(ӊr&        �8�������s�������{���o ?�������ÿ�w�           AD      0 �   `            �               0              @   0 �   `   �������������������?>?�0~G�����|�?ǁ�~>��������>�8�������������������                                                                                                 q�����ߌ9����{�8������ ?��������?��                    0 �   `            �              0               �   0 �   `   ������������������~�����O����������������������������9���?����������������                                                                                                 ���Ï���88�q���w������Ç� � {c���?                     0 �   `          �               0              �   0 �   `   �����������������������������������������������������������?����������������                                                                                                 �8�Ý���8s���wϜ�s��� n �< ����w                     0 �   `         0 �           @   0            �   0 �   `   ������������������������������������������������������������?����������������                                                                                                 q�����π8?8 ��s�8~s��� | �� �����                     0 �   `     @   0 �   `      �   0 �   `     �   0 �   `   ���������������������������������������?�������������������?����������������                                                                                                  ��  ` 00 0    q�8 `    0          �                      0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                      �       0        `                                      ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                <x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       >      <   qς �                                          �����                                                                                                                                                                                                                                                              B   "�(   �                                        (��                                                                                                                                                                                                                                                             @   �(                                             (��                                                                                                                                                                                                                                                        �9$�p @sĴ���/Ă'<z*�                                    9��A(��rb]�9�p                                                                                                                                                                                                                                                <�E$� @�$�P�(�$�Ȣ"�+                                     E$�/�t��RQ(�"                                                                                                                                                                                                               @                                 �}T��0@�$�P� �$�(� ��*                      @              }$�(���BRQ=(" x                                               @                                                                                                                                                                                               �AU� @�$�P� �$�(� ��*                                    A%(��n"RQE(2 �                                                                                                                                                                                                                                              �D�� B�#%P �(�#(���j                                     E%(��2��QE(�"�                                                                                                                                                                                                                                                �8��p <s�$�H>q���<y�                                     9$�A���� a^<��x                                                                                                                                                                                        �                                                                          �                                              �                              �                                                                                                                                                                                                                             �          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             @                                                                               @                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         @                                                                               @                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �                          �                                                   �                          0                                                   �                          0                                                                              �                                                                              ��                 �                                                                             �                                                                             �                                                            ��                                                                             �                                                                             @                                                                            @                                                                           ���                                                                             �                                                                                                                                                                                                                                          ���                                                                            ���                                                                                                                                                                                                                                          ���                                                                            ���                                                                                                                                                                                                                                            ?���                                                                           ���                                                                                                                                                                                                                                     ���                                                                         ���                                                                                                                                                                                                                                    ����                                                                           ���                                                                                                                                                                                                                                    ����                                                                       �    ���                                     �                                 �                                            �                                 �                                            �                                     �����                                                                           ����                                                                            �                                                                            �                                                                        �����                                                                          ���                                                                              �                                                                              �                                                                         �����                                     �                                   '���                                      �                                     �                                      �                                     �                                                                         �����                                                                           ���                                                                              �                                                                              �                                                                         �����                                                                           ���                                                                              �                                                                              �                                                                         �����                                                                          @���                                                                             �                                                                             �                                                                         �����                                                                         ���                                                                             �                                                                             �                                                                         �����                                                                           ��                                                                               �                                                                               �                                                                         �����                                                                         ��                                                                              @                                                                              @                                                                         �����                                                                          /N��                                                                               �                                                                               �                                                                         �����                                                                         /� ?�                                                                              �                                                                              �                                                                         �����                                                                        o���                                                                             �                                                                             �                                                                         �����                                                                         ����                                                                              0                                                                              0                                                                         �����                                                                         ?N��                                                                             �                                                                             �                                                                        �����                                                                         ��                                                                            0                                                                            0                                                                        �����                                                                         ��                                                                              �                                                                              �                                                                         �����                                                                         	����                                                                              `�                                                                              `�                                                                         �����                                                                         ����                                                                              ��                                                                              ��                                                                         �����                                                                         I����                                                                            ��                                                                            ��                                                                         �����                                                                         ����                                                                           ��                                                                           ��                                                                        �����                                                                         ����                                                                            �                                                                            �                                                                         �����                                                                         ���                                                                           � �                                                                           � �                                                                          �����                                                                          �?��                                                                            � ?�                                                                            � ?�                                                                          ����                                                                           ���                                                                            ���                                                                            ���                                                                           ����                                                                           ?���                                                                            ;���                                                                            ;���                                                                           ���                                                                           ���                                                                            ���                                                                            ���                                                                           ?���                                                                           ���                                                                            ���                                                                            ���                                                                           ���                                                                           ���                                                                            ���                                                                            ���                                                                           ���                                                                           ���                                                                            ���                                                                            ���                                                                           ���                                                                            ��                                                                             ��                                                                             ��                                                                             ��                                                                             �                                                                              ?�                                                                              ?�                                                                             �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                     ��                       @                                                     ��                       @                                                                                                                                                                                                           @         ��                       @                                           @         ��                       @                                                                                                                                                                                                           @         ��                       @                                           @         ��                       @                                                                                                                                                                                                           @         ��                       @                                           @         ��                       @                                                                                                                                                                                                           @         ��                     ����                                         @         ��                     ����                                                                                                                                                                                                         @         ��                     ����                                         @         ��                     ����                                                                                                                                                                                                         @         ��                     ?����                                         @         ��                     ?����                                                                                                                                                                ���������                               @         ��                     �������������                               @         ��                     ����                                                                                                                                                                ���������                               @         ��                     ��������������                               @         ��                     �����                                                                                                                                                                ���������                      |         @         ��                    ��������������                      |         @         ��                    �����                                                                                                                                                                ���������                      |         @         ��                    ��������������                      |         @         ��                    �����                                                                                                                                                                ���������                      |         @        ��                    ��������������                      |         @        ��                    �����                                                                                                                                                                ���������                      �         @        ��                    ��������������                      �         @        ��                    �����                                                                                                                                                                ���������                      �      �������     ��                    ��������������                      �      �������     ��                    �����                                                                                                                                                                ���������                      �      �������     ��                    ?��������������                      �      �������     ��                    ?�����                                                                                                                                                                ����������                    �      �������     ��                    ���������������                    �      �������     ��                    �����                                                                                                                                                                ����������                    �      �������     ��                    ����������������                    �      �������     ��                    ������                                                                                                                                                                ����������                    �     �������     ��                   ����������������                    �     �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ?����������������                    ��    �������     ��                   ?������                                                                                                                                                                �����������                   ��    �������     ��                   �����������������                   ��    �������     ��                   ������                                                                                                                                                                �����������                   ��    �������     ��                   ������������������                   ��    �������     ��                   �������                                                                                                                                                                �����������                   ��    �������     ��                  ������������������                   ��    �������     ��                  �������                                                                                                                                                                �����������                   ��    �������     ��                  ������������������                   ��    �������     ��                  �������                                                                                                                                                                �����������                  ��    �������     ��                  ������������������                  ��    �������     ��                  �������                                                                                                                                                                �����������                  ��    �������     ��                  ������������������                  ��    �������     ��                  �������                                                                                                                                                                �����������                  ��    �������     ?��                  ������������������                  ��    �������     ?��                  �������                                                                                                                                                                �����������                  ��    �������     ?��                  ������������������                  ��    �������     ?��                  �������                                                                                                                                                                ������������                  ��    �������     ?��                  �������������������                  ��    �������     ?��                  �������                                                                                                                                                                ������������                  ��    �������     ?��                  �������������������                  ��    �������     ?��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            