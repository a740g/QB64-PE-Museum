�P  �6>+ ����������������������������������������                                        ����������������������������������������                                        �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ��������������������������  >  |   ����                                                                               �                          ���������   ������������������������������}��������                          ���������                              ��������   �  �    ��0 �  �      � ���������   ������������������������������}��������  �    ��0 �  �      � ���������      �    ��0 �  �      � ��������   �      �0 �0 �      ` ���������   ������������������������������}��������      �0 �0 �      ` ���������          �0 �0 �      ` ��������   �      �0 �0 �      ` ���������   ������������������������������}��������      �0 �0 �      ` ���������          �0 �0 �      ` ��������   �  �y������9����>͛6l ���������   ������������������������������}��������  �y������9����>͛6l ���������      �y������9����>͛6l ��������   �  �l̀0ͳ;��0Ͷ�3f͛6` ���������   ������������������������������}��������  �l̀0ͳ;��0Ͷ�3f͛6` ���������      �l̀0ͳ;��0Ͷ�3f͛6` ��������   �  l���ͳ3ϳ�Ͷ۳f�͛6` ���������   ������������������������������}��������  l���ͳ3ϳ�Ͷ۳f�͛6` ���������      l���ͳ3ϳ�Ͷ۳f�͛6` ��������   �  l��0ͳ3ٳ Ͷ�3f͛6` ���������   ������������������������������}��������  l��0ͳ3ٳ Ͷ�3f͛6` ���������      l��0ͳ3ٳ Ͷ�3f͛6` ��������   �  l̓0ͳ3ٳ0Ͷ�3f�` ���������   ������������������������������}��������  l̓0ͳ3ٳ0Ͷ�3f�` ���������      l̓0ͳ3ٳ0Ͷ�3f�` ��������   �  �fy�����ϙ�Ͷ�>l ���������   ������������������������������}��������  �fy�����ϙ�Ͷ�>l ���������      �fy�����ϙ�Ͷ�>l ��������   �               �    ` ���������   ������������������������������}��������               �    ` ���������                   �    ` ��������   �               �    8p� ���������   ������������������������������}��������               �    8p� ���������                   �    8p� ��������   �                          ���������   ������������������������������}��������                          ���������                              ��������   �                          ���������   ��������������������������  >  |   ����                          ���������                                           �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                                                               �                                                                                                                                               ?��� ���������������  ?  ��������� �  ����?���>+ ����������������������������������������                                        ����������������������������������������                                        �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ��������������������������  >  |   ����                                                                               �                          ���������   ������������������������������}��������                          ���������                              ��������   �  ?              0`    ���������   ������������������������������}��������  ?              0`    ���������      ?              0`    ��������   �  0 �     `    0`    ���������   ������������������������������}��������  0 �     `    0`    ���������      0 �     `    0`    ��������   �  0 �     `    0`    ���������   ������������������������������}��������  0 �     `    0`    ���������      0 �     `    0`    ��������   �  0|�yϞp|����lٳf����������   ������������������������������}��������  0|�yϞp|����lٳf����������      0|�yϞp|����lٳf���������   �  >v����`�3�m�6`lٳf ���������   ������������������������������}��������  >v����`�3�m�6`lٳf ���������      >v����`�3�m�6`lٳf ��������   �  0f��}��`��?�m�6nlٳf ���������   ������������������������������}��������  0f��}��`��?�m�6nlٳf ���������      0f��}��`��?�m�6nlٳf ��������   �  0f�3͙�`͛0�m�6`lٳf ���������   ������������������������������}��������  0f�3͙�`͛0�m�6`lٳf ���������      0f�3͙�`͛0�m�6`lٳf ��������   �  0f��3͙�`͛3�m�6`8p�� ���������   ������������������������������}��������  0f��3͙�`͛3�m�6`8p�� ���������      0f��3͙�`͛3�m�6`8p�� ��������   �  ?fg�}��0|���m���0`������������   ������������������������������}��������  ?fg�}��0|���m���0`������������      ?fg�}��0|���m���0`�����������   �         �         0`�� ���������   ������������������������������}��������         �         0`�� ���������             �         0`�� ��������   �                   �Ç ���������   ������������������������������}��������                   �Ç ���������                       �Ç ��������   �                          ���������   ������������������������������}��������                          ���������                              ��������   �                          ���������   ��������������������������  >  |   ����                          ���������                                           �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                            `      ~����             �       �                                       ����������������������������������������                                            0` `    `�1�`   �       �0      �                                       ����������������������������������������                                            0` `    `�1�`   �       �0      �                                       ����������������������������������������                                            0l�p��p`�1�s����<�����9�      �                                       ����������������������������������������                                            0l�`͙��|�1��fa���٘f͙����3      �                                       ����������������������������������������                                            0l�`͟�``�1�fa�����`͙�6ϳ�      �                                       ����������������������������������������                                            3l�`͘0`�1�fa��ـ`͙�6ٳ      �                                       ����������������������������������������                                            3m�`͙��`�1�fa���٘fݙ�6ٳ3      �                                       ����������������������������������������                                            1��0��p~�1�3��g��<}��3ϙ�      �                                       ����������������������������������������                                            0   �                             �                                       ����������������������������������������                                               �                             �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                       ����������������������������������������                                                                               �                                                                               �                                                                                                                                                                                                   