�P   N � ���������������������������������������������������������������������������������������������������������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �?������������������������������?����������������������������� ��                            ������������������������������� �                             �                              ��                            ��                             �/������������������������������/����������������������������� ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                        ����(�(                        ����( ��                        ����������������������������������� �(                        ����(�(                        ����( ��                        ��������������������������������� �( �9��O>�Bp              ����(�( �9��O>�Bp              ����( �� �9��O>�Bp              �����������������������������?�� �( �DD(P��b�              ����(�( �DD(P��b�              ����( �� �DD(P��b�              �?���������������������������� �� �( �@D(P�b�              ����(�( �@D(P�b�              ����( �� �@D(P�b�              � �������������������������������� �( �@D(P�R�              ����(�( �@D(P�R�              ����( �� �@D(P�R�              ����������������������������������� �(                        ����(�(                        ����( �� �8G�P�Rp              ����������������������������������� �(                           (�(                           ( �� �D(P�J              ������������������������������� �� �(                         �� (�(                         �� ( �� �D(P�F              � ����������������������������?�� �(                        �� (�(                        �� ( �� �DD(P��F�              �?������������������������������ �(                        �� (�(                        �� ( �� �8D'��Bp              ��������������������������������� �(                            (�(                            ( ��                        ����������������������������������� �(                            (�(                            ( ��                        ����������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( �� �           
     @     ���w������������������������� �(                            (�(                            ( �� �    �          @�   ���w������������������������� �(                            (�(                            ( �� �    �         @�   ���v?��?1�i�~S��������}�1���� �(                            (�(                            ( �� ��dY���8䁬p��sg$�x��v  ����k��n������w������[}��n���� �(                            (�(                            ( �� � �R �YE2�� 
H��E�I  ���t��n�����������U}��n���� �(                            (�(                            ( �� ��DS��}"�
�� zH��E�I  ���u�ۭ�n���������u�U}��n���� �(                            (�(                            ( �� � $R �A"�
�� �H��E�I  ���u�k-�n����~�w����u�n���n���� �(                            (�(                            ( �� � �� �QE�"�B� �H�E�I  ���?��?��n��]��������������� �(                            (�(                            ( �� ��cQ�N�8�@�pB��zGx�NI  ������������������������������� �(                            (�(                            ( ��                           ������������������������������� �(                            (�(                            ( ��                           ������������������������������� �(                            (�(                            ( ��                            ����������������������������� �(                            (�(                            ( ��      @       @        @ ���������~��������������������� �(                            (�(                            ( ��      �      @        @���������~��������������������� �(                            (�(                            ( ��      �      @        @�����4�g�>S���4����Lm�4�m��O� �(                            (�(                            ( �� q�3���p�q�X�9��@��`x����u�[��~�w��u�o����ۭ��]mo��7� �(                            (�(                            ( �� �,�P"�2�%�,�e$RA,���E����|X/�~���o���۪�w]U���w� �(                            (�(                            ( �� ���"�"���E�=$U@���@E����}�[��~���}�o����۪��]Uߺ�w� �(                            (�(                            ( �� ��"�"�	��E E$U@H�� E����u�[��~�w��u�o���۷~�]�o��w� �(                            (�(                            ( �� �(�P"�"�%�(�EE$H�(�D�E�����7lo�]���7k����w7c���w� �(                            (�(                            ( �� qȓ���p�qȔD�=#��ȜD`x�������������������������������� �(                            (�(                            ( ��                           ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��  @            !   ���o�������������������������� �(                            (�(                            ( �� �           $ 	    I   ���o�������������������������� �(                            (�(                            ( �� �           $ 	    I   ���)��8�p�ɍ8J�~ڧ���� �(                            (�(                            ( �� �8Y�4��6rǵ��c�%X�Mc� ���f���Z���[t�Y���k�ښ�k��� �(                            (�(                            ( �� �DR(�@Q��(�A	�A%eI�@ ���n��������[����>����?�� �(                            (�(                            ( �� �|S�%@�Q$�(�A	�UEI� ���n��������}�[������������ �(                            (�(                            ( �� �@R%AQ$�(�A	UEI  ���n���Z���[u�[����v����� �(                            (�(                            ( �� �DR(�AQ��(�A	@�EI@ ������8������k���v����� �(                            (�(                            ( �� Q8Q��@�Or'�@���D�E� ������������������������������ �(                            (�(                            ( ��               �        @   ������������������������������� �(                            (�(                            ( ��                           ������������������������������� �(                            (�(                            ( ��                            ����������������������������� �(                            (�(                            ( �� �         �         P  ����������������������������� �(                            (�(                            ( �� �   H     �     $    H  ���������������������������� �(                            (�(                            ( �� �   H     �     $    H� ���cNϔ��ɍ��N?�1�g�q�j�7��� �(                            (�(                            ( �� ���0k6rH��f�X�5��c�� ���]5�_�]�[u��5�kn��ٮ�jk����� �(                            (�(                            ( �� ��(�L� ��H� ��eP&Q��H@ ���]u�_�A�[uW�t�n��/۠������� �(                            (�(                            ( �� ��/�H������D�E�$_UH@ ���]u�߷_�[uW�u��n���ۯ����?�� �(                            (�(                            ( �� ��( H����� $�E$PUH� ���]u�_�]�[v��u�kn��ۮ������� �(                            (�(                            ( �� ��(�H���� ��EP$Q%H  ���cv��c�[���v?�q�o����5���� �(                            (�(                            ( �� ��� (��q��b�D�N%�  ������������������������������� �(                            (�(                            ( ��                         �����?������������������������ �(                            (�(                            ( ��  �            �         ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( ��           �       A    ������������������������������� �(                            (�(                            ( ��                  A    ������������������������������� �(                            (�(                            ( ��                  A    ����1��q�NmS��?�2�ko����8�� �(                            (�(                            ( �� f�X�9�2����xr�q���y9$� ���kn��뮵5�mMw������o������ �(                            (�(                            ( �� ��eEQJ� ���" 
)T�EE$(�����n����u�U]w߅߅��+o������ �(                            (�(                            ( �� D�EEQ"� ��� z z	ԐEET/�����n����u�U]w�u�u��o������� �(                            (�(                            ( �� $�EEQ� ��� � �	T�EET( ���kn��뮵u߻]w�u�u�˫���w��� �(                            (�(                            ( �� ��EEQJ� D��"� �)4T`ED�(�����q��q�v�]��߆;,+���w���� �(                            (�(                            ( �� b�D�9�2��D�xz y���@y8�
' ������������������������������� �(                            (�(                            ( ��                  @      �����������?����������������� �(                            (�(                            ( ��   �  �         �      ������������������������������� �(                            (�(                            ( ��                            �������������o�������������� �(                            (�(                            ( �� �    �     � �         �������������߷�������o������ �(                            (�(                            ( �� �    �      H     @�    �������������߷�������o������ �(                            (�(                            ( �� �    �      H     @�    ���4�N?8�m��?O����1��)��9��� �(                            (�(                            ( �� ������$�s<��k�8`�8�0 ���w�}7�w�Wm���_�]��n��f��ַ�� �(                            (�(                            ( �� �,�� �(��
E �L�"�D@�D)H ���vavv�U��_�A��o��n������ �(                            (�(                            ( �� �螉���0�zD��H�"�|@�|$  ���u�]u�u��Uu��_�_��o��n������ �(                            (�(                            ( �� �(�� �((��D@�H�"�@@�@" ���u�]u�u�[�u��_�]��n��n��ַ�� �(                            (�(                            ( �� �(�� �(�D�E �H�"�D@�D)H ���avݻ��?_�c��q����9��� �(                            (�(                            ( �� �螉���"Dz<��(��8@Q8	�0 ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( �� �                       ������������������������������� �(                            (�(                            ( ��                        ������������������������������� �(                            (�(                            ( ��                        ���f�~dƜ?q�
o���������������� �(                            (�(                            ( �� �a��9c��D��               ���Zn���k�鮺����������������� �(                            (�(                            ( �� ��RE�AQEP               ���n����������������������� �(                            (�(                            ( �� �EA�QEP               ���v��m���������������������� �(                            (�(                            ( �� � �EAQEP               ���Z�����뮲����������������� �(                            (�(                            ( �� �REAQM@               ���f�~u��?������������������� �(                            (�(                            ( �� ���9��N4�P               ������������������������������� �(                            (�(                            ( ��       @                   ����������������������������� �(                            (�(                            ( ��      �  �                ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                 � @ @   (�(                 � @ @   ( ��                 � @ @   ������������������������������� �(                 @ @ @   (�(                 @ @ @   ( ��                 @ @ @   ������������������������������� �(                   @ @   (�(                   @ @   ( ��                   @ @   ������������������������������� �(                 8�A�@   (�(                 8�A�@   ( ��                 8�A�@   ������������������������������� �(                 	�EAT@   (�(                 	�EAT@   ( ��                 	�EAT@   ������������������������������� �(                 QEA@   (�(                 QEA@   ( ��                 QEA@   ������������������������������� �(                 QEA@   (�(                 QEA@   ( ��                 QEA@   ������������������������������� �(                 �EA4R    (�(                 �EA4R    ( ��                 �EA4R    ������������������������������� �(                 N8�|ӑ@   (�(                 N8�|ӑ@   ( ��                 N8�|ӑ@   ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ��                             �/������������������������������/����������������������������� ��                            ������������������������������� �                             �                              ��                            ��                               �?������������������������������?����������������������������� ��                            ��                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ��������������������������������                                ��������������������������������                                ��������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            