�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?����������������������������������������������������o���W����������������������������o���W����������������������������o���W���������?�����������������������������������{������������ۿ������������������{������������ۿ������������������{������������ۿ����������������?�����������������������������������������������ۿ������������������������������ۿ������������������������������ۿ����������������?�����������������������������������1��Lm�p��q�4�۱��鍏��9����������1��Lm�p��q�4�۱��鍏��9����������1��Lm�p��q�4�۱��鍏��9��������?�����������������������������������~�~��_����鮵�[�n���uw��ֻ���������~�~��_����鮵�[�n���uw��ֻ���������~�~��_����鮵�[�n���uw��ֻ�������?�����������������������������������~p��\*���믵�oۮ���}��ۃ���������~p��\*���믵�oۮ���}��ۃ���������~p��\*���믵�oۮ���}��ۃ�������?�����������������������������������~�n��[����믵�wۮ���}��ݿ���������~�n��[����믵�wۮ���}��ݿ���������~�n��[����믵�wۮ���}��ݿ�������?�����������������������������������z�n��[�k��ˮ��[ۮ���uw��ֻ���������z�n��[�k��ˮ��[ۮ���uw��ֻ���������z�n��[�k��ˮ��[ۮ���uw��ֻ�������?���������������������������������������\7k��+��7g�q��k���T9�������������\7k��+��7g�q��k���T9�������������\7k��+��7g�q��k���T9�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������}����������������������������������}����������������������������������}��������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������}N?p����Ɵ�6�}����>Q8��������}N?p����Ɵ�6�}����>Q8��������}N?p����Ɵ�6�}����>Q8������?�����������������������������������}5���_Z���ot���ֺ���ku���[�������}5���_Z���ot���ֺ���ku���[�������}5���_Z���ot���ֺ���ku���[�����?�����������������������������������}t��Xn}���u���=ۂ�����o�������}t��Xn}���u���=ۂ�����o�������}t��Xn}���u���=ۂ�����o�����?�����������������������������������}u����v���u����ݾ�u��}�����������}u����v���u����ݾ�u��}�����������}u����v���u����ݾ�u��}���������?�����������������������������������}u����Z���u�>뽖��u��u���[�������}u����Z���u�>뽖��u��u���[�������}u����Z���u�>뽖��u��u���[�����?�����������������������������������v?���f�����~~Y����?V���������v?���f�����~~Y����?V���������v?���f�����~~Y����?V�������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?��������������������������������������cO��yN9��3cN���������������cO��yN9��3cN���������������cO��yN9��3cN����������?�����������������������������������m��V��]7��5ֻ�u��]5��]����������m��V��]7��5ֻ�u��]5��]����������m��V��]7��5ֻ�u��]5��]��������?�����������������������������������m��V�]w��t��t]v��Aꮳ���������m��V�]w��t��t]v��Aꮳ���������m��V�]w��t��t]v��Aꮳ�������?�����������������������������������mu�V��]w��u���u��]w�_ꮵ���������mu�V��]w��u���u��]w�_ꮵ���������mu�V��]w��u���u��]w�_ꮵ�������?�����������������������������������mu�V��]w��uֻ�u��]u��]�n����������mu�V��]w��uֻ�u��]u��]�n����������mu�V��]w��uֻ�u��]u��]�n��������?�����������������������������������m�V�cu���v9��7cvw�c�q���������m�V�cu���v9��7cvw�c�q���������m�V�cu���v9��7cvw�c�q�������?���������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������?���������������������������������?���������������������������������?�����������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������W�������������������������������W�������������������������������W�������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������mW͵1��t�'c�m�>Sg�p�p�����������mW͵1��t�'c�m�>Sg�p�p�����������mW͵1��t�'c�m�>Sg�p�p�������?��������������������������������������mW��n��u���]�m���[ۮ��������������mW��n��u���]�m���[ۮ��������������mW��n��u���]�m���[ۮ���������?�������������������������������������UW�Uo��u��_�m���o�.��.�����������UW�Uo��u��_�m���o�.��.�����������UW�Uo��u��_�m���o�.��.�������?�����������������������������������u��UW�Uo��u���_um���w�������������u��UW�Uo��u���_um���w�������������u��UW�Uo��u���_um���w�����������?�����������������������������������u��W��n��e���]us���[ۮ�����������u��W��n��e���]us���[ۮ�����������u��W��n��e���]us���[ۮ���������?��������������������������������������W�����c�w�?]g�p�p������������W�����c�w�?]g�p�p������������W�����c�w�?]g�p�p�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�������������������������������������jq��q�og�f8�������������������jq��q�og�f8�������������������jq��q�og�f8���������������?�����������������������������������k�{i��ٮ��[���������������������k�{i��ٮ��[���������������������k�{i��ٮ��[�������������������?�������������������������������������z���۠��o�
��������������������z���۠��o�
��������������������z���۠��o�
����������������?������������������������������������w����ۯ��w�����������������������w����ۯ��w�����������������������w����ۯ��w��������������������?�����������������������������������j�}ۮ�ۮ��[���������������������j�}ۮ�ۮ��[���������������������j�}ۮ�ۮ��[�������������������?�������������������������������������۱���og�v8_�������������������۱���og�v8_�������������������۱���og�v8_���������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������{~������������������������������{~������������������������������{~����������������������������?�����������������������������������:�w������������������������������:�w������������������������������:�w����������������������������?�����������������������������������:�w�w���������������������������:�w�w���������������������������:�w�w�������������������������?�����������������������������������Z�w�wq���8��e���8cm�S��1���������Z�w�wq���8��e���8cm�S��1���������Z�w�wq���8��e���8cm�S��1�������?�����������������������������������Z�p�w~�M��{_�����]m���w��n��_������Z�p�w~�M��{_�����]m���w��n��_������Z�p�w~�M��{_�����]m���w��n��_����?�����������������������������������j�w������}�-��U�]U����n��_������j�w������}�-��U�]U����n��_������j�w������}�-��U�]U����n��_����?�����������������������������������r�w�������ۭ��U�]U����n��_������r�w�������ۭ��U�]U����n��_������r�w�������ۭ��U�]U����n��_����?�����������������������������������r�w���]��{[�����]���w��n��_������r�w���]��{[�����]���w��n��_������r�w���]��{[�����]���w��n��_����?�����������������������������������{p_��������6Y���c���]������������{p_��������6Y���c���]������������{p_��������6Y���c���]����������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������o���������������������������������o���������������������������������o�������������������������������?�����������������������������������o���������������������������������o���������������������������������o�������������������������������?�����������������������������������)���4���|���~8�&7��9�P��������)���4���|���~8�&7��9�P��������)���4���|���~8�&7��9�P������?�����������������������������������f���u�{u�k�����Mm�ouֺ�Z��������f���u�{u�k�����Mm�ouֺ�Z��������f���u�{u�k�����Mm�ouֺ�Z������?�����������������������������������n���{u��=��v��]m׿t��Z��������n���{u��=��v��]m׿t��Z��������n���{u��=��v��]m׿t��Z������?�����������������������������������n���}�{u�����v��]m��u���Z��������n���}�{u�����v��]m��u���Z��������n���}�{u�����v��]m��u���Z������?�����������������������������������n���u�{u�뽺��˽�]m�ouֺ�Z��������n���u�{u�뽺��˽�]m�ouֺ�Z��������n���u�{u�뽺��˽�]m�ouֺ�Z������?���������������������������������������7{���~��+�8ݮ7��9���������������7{���~��+�8ݮ7��9���������������7{���~��+�8ݮ7��9���������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        