�P  X�/ / ��� � p�������  �  ���  3��������  �  ��Ç�F ������Ç��  ?�  �����������~������  ?�  ����i�������������  ?�  ��Ài���Ç����Ç��  ?�  ���o�� ��N�����  �  � 7�� ���� � ��� ����^���?�����?� ��� ����� � ����  � ��� ���7��`�?~��  ?� ��� ����� t���  � ��� ������t���  � ��� E�;���:����  �� ��  �^E����:����  �� ��  �x"�7������� ��  ��  � �������2����� ��  ����}� �  ���  � ��� ����< ��������?� ��� ������ ����������� ��� ����?����� �����?� ��� ����    ~��  � ��� �������   >�����  ?�  �������   6�����  ?�  ���g��� � �����  ?�  ���3��p �  �����  �  ���3��  �  �����  �  ���3��  �? �����  �  �����  �?������  �  ��>��  ?�?���>��  ��  ��>��  ?����>��  ��  ��?��  ?����?��  ��  ��?���     �� ��  ��  ��~��  �� ��~ �� ��  ��������  ����� ��� �y��?����� ����?� ��� �y�?�����  ��� ?� ��� �3������� ��� � ��� �������� ��� � ��� ���������� � ��� ���?��������� � ��� � ��?���L��  � ��� �������   ��  � ?���  ��������� ������ ?��� @�������0 ��� � ?��� ��������0 ��� � ?��� l�������0 ��� � ?���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ���pi�����������  �  ��o�� ��N�����  �  � �������� �� ��  ����W^��������� ��� ���k����������c�� ��� ��w�7��`��?~��s�?� ��� ����� t���  � ��� ������t���  � ��� E�;���:����  �� ��  �^E����:����  �� ��  �x"�7������� ��  ��  � �������2����� ��  ����}� �  ���  � ��� ����< ��������?� ��� ������ ����������� ��� ����?����� �����?� ��� ����    ~��  � ��� �������   >�����  ?�  �������   6�����  ?�  ���g��� � �����  ?�  ���3��p �  �����  �  ���3��  �  �����  �  ���3��  �? �����  �  �����  �?������  �  ��>��  ?�?���>��  ��  ��>��  ?����>��  ��  ��?��  ?����?��  ��  ��?���     �� ��  ��  ��~��  �� ��~ �� ��  ��������  ����� ��� �y��?����� ����?� ��� �y�?�����  ��� ?� ��� �3������� ��� � ��� �������� ��� � ��� ���������� � ��� ���?��������� � ��� � ��?���L��  � ��� �������   ��  � ?���  ��������� ������ ?��� @�������0 ��� � ?��� ��������0 ��� � ?��� l�������0 ��� � ?��� ������            �����������            �����~������            �����~������            �����>������            �����>������            ������������            �����������            ����������            #��������            ��o?������            9�����?����            ����������            �����������            ���� �����            ��������?��  / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ���׀�X �������  �  ������c��~�����  �  ��ϟ�� � �������  �  ������Ã���������  ?�  ��;���G���������  ?�  �_���������������  ?�  �x9�7�������������  �  � <��������2������  �  ���K�� �<s����C��  �  ���� �>s������  �  ��ޗ�� �g������  ?�  ���1����� ������  ?�  ������  ~�����  �  �������   >�����  �  �������   6�����  �  ������ � �����  ��  ����p �  ���� ��� ����?�      ��  ?� ��� ����� ��� ����� ��� ��� =�  ��?���� ?� ��� ����    ?���  � ��� ������   ������  �  ������   ������  �  ���7��  �  �����  �  �����  �� �����  �  �������� �����  ?�  ���������������  �  �������  � �����  �  �??����?�� ��? ��  ��  ������  ���� ��� ����?� �� ����?� ��� ���?�������� ?� ��� ��??�?������ ?� ��� ��������  ��� � ���  ������    ��  � ��� @��������� ������ ��� ��������  ��� � ��� l�������  ��� � ��� ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      ������Á@��������      ��;��� ��������      �_���������������      �x�7���� ��������      � ������p�2������      ������ �?��������      ����� �8��������      ������ � �������      ��������  �������/ / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      �?�����@����?��� �   ��;���� �������� �   �\�?���| ����\?�� ��  �y��7����������� ��  ����������2������ ��  ������ ��{����{�� ��  ��=� �������� ��  ��?��� ������?��� ��  �������� ����� ��� ������ ~���� ��� ����?���� >����?� ?��� ����?���� 6����?� ?��� Ϗ����?�������� ��� �����p=��� ����� ��� �?���� ~��� �>��� ���� �]���� O�� �M�� ���� �p7�� C��@�� ���� ��O�?� ?�?����?� ��� �ȟ�� ������ ?��� ��~�  �����~� ��� ����� ��  ����� ��� ������ ��� ������ ��� ������    ��  � ��� �s��?����� ����?� ��� �y�����  @ ��  � ��� �> 9������ �� �� ��  ��������  ����� ��  ������� ��� �� ��  ������������ �� ��  ���?������ � ��� ���?����  �� ?� ���  ������    ��  ?� ��� @��������� ������ ��� ��?������@ ��� � ��� l�?������@ ��� � ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      �0��   ���0� �� �7���������7�� �� 7�;��������7�� �� �]���������7�� �� �y�7���������� ��� ��w�����2���� ��� ���}� �������� ��� ���| �������� ��� ���� �������� ��� �������� ����� ��� �����    ~��  � ��� ��?����   >�� ��  ��  �������   6�����  ?�  �������   �����  �  �����p �  �����  ��  ��  ��  ��  ��  �� ��  ����}� ��? ����� ��� �����    ?���  �� ��  ������    ?������  �  ������   ������  �  �����  �������  �  ������  �  ������  �  �����  �� �����  �  ��������� ������  ?�  ���������������  ?�  �������  � �����  ?�  �?�����?� �����  �  �������  �����  ��  ������ �� ������ ��  ������������ �� ��  ��>��?������ �� ��  �������  ��� � ���  �����    ��  � ��� @��������� ������ ��� ��������  ��� � ��� l�������  ��� � ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      ������Á@��������      ��;��� ��������      �_���������������      �x�7���� ��������      � ������p�2������      ������ �?��������      ����� �8��������      ���g�� � ������  �  ��������� �������  �  ������ � ~������  �  ������� � >������  �  ������� � 6������  �  ������� � ������  �  �����p �  �����  �  �����  �  �����  �  ���?��  �? ���?��  �  ������   ?����?��  �  ������    ?������  ?�  ������  ?��������  �  ��Ç��   ������  ?�  ������   3  ���?��  �  ������  �� ������  �  �������� �����  �  �������������  �  �������  � �����  ?�  �?�����?� �����  �  �������  �����  ��  ������ �� ������ ��  ������������ �� ��  ��?�?������ � ��� �������  ��� � ���  �����    ��  � ��� @��������� ������ ��� ��������  ��� ?� ��� l�������  ��� ?� ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  <p�������  �  ���?�F �<t�������  �  ���������~�����  �  ���i�����������  �  ���pi�����������  �  ��qo�� �O�N�����  �  ��?���
�����?��  �  ��� �^�� ����`�� ��  ��  W��   ���  � ��� ��  w��`  ~��  � ��� �  ���   ����  �� ��  � ����  ���� �� ��   ;���  ���� ��  ��  �_����� �������  �  �x 7���� �������  �  �  ����  �2�� ��  ��  ��| �� �| ���c��� ��  ��  | �  ���  � ��� ��� ?� �� �����?� ��� ��  ���   ���  � ��� ��	���   ~�����  �  ������   >�����  �  ������   6�����  �  ������   �����  �  �����p    �����  ?�  �����     �����  ?�  �����   ? �����  ?�  �����   ?������  ?�  �����    ?������  �  �����   ������  �  �����   ������  �  �����     �����  �  ��<��  < � ��#���  ��  ��x ���x � ��t�� ��  �|� ����  ���� ��� �|� ���� @ ��H �� ��� �<` ���`   ��� �� ��� ��  ��    ��  �� ��� ��  ?�    ��  � ��� ��  ?��  ���  � ��� �   �?�  ��  ?� ��� �� ����  ���� ���     ���    ��  � ��� @   ���    ��  � ��� �   ���    ��  � ��� l   ���    ��  � ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� �O�N�����  �  ��?���
�����?��  �  ��� �^�� �����f�� ��  ��  W��   ����� ��� ��  w��`  ~��  � ��� �  ���   ����  �� ��  � ����  ���� �� ��   ;���  ���� ��  ��  �_����� �������  �  �x 7���� �������  �  �  ����  �2�� ��  ��  ��| �� �| ���c��� ��  ��  | �  ���  � ��� ��� ?� �� �����?� ��� ��  ���   ���  � ��� ��	���   ~�����  �  ������   >�����  �  ������   6�����  �  ������   �����  �  �����p    �����  ?�  �����     �����  ?�  �����   ? �����  ?�  �����   ?������  ?�  �����    ?������  �  �����   ������  �  �����   ������  �  �����     �����  �  ��<��  < � ��#���  ��  ��x ���x � ��t�� ��  �|� ����  ���� ��� �|� ���� @ ��H �� ��� �<` ���`   ��� �� ��� ��  ��    ��  �� ��� ��  ?�    ��  � ��� ��  ?��  ���  ?� ��� �   �?�  ��  ?� ��� �� ����  ���� ���     ���    ��  � ��� @   ���    ��  � ��� �   ���    ��  � ��� l   ���    ��  � ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ���׀�Z ��������  �  ������c�C�~�����  �  ��?��� � �����?��  �  �����Ã ��������  �  �;���b ��������  �  �_����� �������  �  �x7���� �������  ;�  � ����� �2�����  =�  ����� �	������  >�  ����� � ����͇��  ?x  ����� � �������  ?�  �������  ������  �  ��	���   ~�����  �  ������   >�����  �  ���?���  ? 6���?��  �  ������   �����  �  ����p   �����  ��  ��  ��      ��  �� ��  ��x }�  x ? ��g�� ��� ��  ��    ?���  �� ��  �����    ?������  �  �����   ������  �  �����   ������  �  �����     �����  �  �����    � �����  �  ������  � �����  ?�  ������  ������  ?�  ������  � �����  ?�  �?������ ������  �  ��0���0  ��(��  ��  ��p �� p  ��|��  ��  ��x ���x ���$�� ��  �  ��?�  ��x�� ��  �   ���   ��  �� ���     ���    ��  �� ��� @� ����   �� ?� ��� �   ���    ��  ?� ��� l   ���    ��  ?� ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      ������Á@��������      ��;��� ��������  `   �_A����A�����A���  �   �x@?7���@ ����0?��  ��  � ������ �2���� ��  �� �� � ����C�� ��  �� � � ��� �� ��  �� �� � ���`�� ��  ��  ����   ������ ��  �� ���  ~��  � ��� ��  ��   >��� ��� ��  ��   6��� ��� ��  ?��   �� ?� ��� ��  ?�p     �� ?� ��� ��  ?�      ���?� ?��� ��  =�   ? ��h?� ?��� ��@ =�    ?���� ?� ?��� ��� �    ?��Ѡ � ?�� ��  �    ���@� ��� ��� ��  � ��� �� ��  ��  �     ��� � ��� ��� ?�  �   ��x �� ��� ��  ��    �� � ��� �|� ����  ����� ��� �~  ����  � ��  �� ��  �?������ ������  �  ��8���8  ��4��  ��  ��x �� x  ��d�� ��  ��p ���p ����� ��  �  ��?�  ��x�� ��  �   ���   ��  �� ���     ���    ��  �� ��� @� ����   �� ?� ��� �   ���    ��  ?� ��� l   ���    ��  ?� ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      ��8����� �������� ��  �8;���� �����>�� ��  �^�8���� �����>�� ��  �x� 7���� �����>�� ��  � � ����� �2����� ��  ��� �� �� ������ ��  ��� � �� ������ ��  ��� �� �� ������ ��  ��� �����  ������ ��  �� ��� �  ~����� ��  �� ���   >�� ��  ��  ������   6�����  ?�  ������   �����  �  �� ��p    �� ��  ��  ��  ��      ��  �� ��  ��� }� � ? ���� ��� ��  ��    ?���  �� ��  �����    ?������  �  �����   ������  �  �����   ������  �  �����     �����  �  �����    � �����  �  ������  � �����  ?�  ������  ������  ?�  ������  � �����  ?�  �?������ ������  �  ��8���8  ��$��  ��  ��x �� x  ��v�� ��  ��x ���x ���&�� ��  �  ��?�  ��x�� ��  �   ���   ��  �� ���     ���    ��  �� ��� @� ����   ��?� ��� �   ���    ��  ?� ��� l   ���    ��  ?� ���                                                                                                                                                                                                                                                                                                                                                                                 / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      ������Á@��������      ��;��� ��������      �_���������������      �x�7���� ��������      � ������p�2������      ������ �?��������      ����� �8��������      ������ � �������      ���q����  ������  �  ��9���  ? ~���?��  �  ������  >�����  �  ������  6������  �  ������  �����  �  �����p    �����  �  �����     ���?��  �  �����   ? �����  �  �����   ?������  �  �����    ?������  ?�  �����  >�������  �  �����   ������  ?�  �����   3  �����  �  ���?��    � ���?��  �  ���?���  � ���?��  �  ������  ������  �  ������  � �����  �  �?������ ������  ?�  ������  �����  �  ��8�� 8  ��>��  ��  ��8���8 �����  ��  � ��?�  ��<��  ��  �   ����   �� �� ��      ����    �� �� ��  @� ?����   ����� ��� �   ?���    ��  � ��� l   ?���    ��  � ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x��� �        �  ��Ï�����  �    �  �Ã���Ç�F  �    ?�  ?|�>�������  �    ?�  |�
����i�  �    ?�  ~��&��Ài�  �    ?�  ��C������o�  �    �  �� H8��7�      ��� }���(�����^ ��   ��� ��~��� ��       ��� ������7�       ��� ����`�t�       ��� �|�� <�t�       ��� ��E��<:;�       ��  �E��|�^:�       ��  0�"��|�x	7�        ��  ���� ���  �   ��  �x��r6��  }�       ��� �y��?�����< ��   ��� �s���|������ ���  ��� ?y��?~����?� ��   ��� �����  �       ��� {����և����        ?�  s����ȏ����        ?�  7��`����χ��        ?�  ���0��������       �  ���0��������       �  ���2��������       �  ����~������       �  ��>�~��?���  >     ��  ��>�>��?���  >     ��  ��?�>��?���  ?     ��  ��?����� ��        ��  ��~������  ~    ��  �|��������  ��   ��� #���?��y��?� ��   ��� ��?��y��?� �    ��� 9����3���� �    ��� �s������� �    ��� ���������� �    ��� ��? ������ �    ��� �� �����O�      ��� ������   '�       ?��� ������ ���� ���  ?��� �����@��7� �    ?��� _�������7� �    ?��� �����l��7� �    ?���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~8�&���pi�        �  ��C�����o�       �  �� H8����      ��  }���(�����W^ ��   ��� ��k�~������ �c�  ��� �w������7�  s�   ��� ����`�t�       ��� �|�� <�t�       ��� ��E��<:;�       ��  �E��|�^:�       ��  0�"��|�x	7�        ��  ���� ���  �   ��  �x��r6��  }�       ��� �y��?�����< ��   ��� �s���|������ ���  ��� ?y��?~����?� ��   ��� �����  �       ��� {����և����        ?�  s����ȏ����        ?�  7��`����χ��        ?�  ���0��������       �  ���0��������       �  ���2��������       �  ����~������       �  ��>�~��?���  >     ��  ��>�>��?���  >     ��  ��?�>��?���  ?     ��  ��?����� ��        ��  ��~������  ~    ��  �|��������  ��   ��� #���?��y��?� ��   ��� ��?��y��?� �    ��� 9����3���� �    ��� �s������� �    ��� ���������� �    ��� ��? ������ �    ��� �� �����O�      ��� ������   '�       ?��� ������ ���� ���  ?��� �����@��7� �    ?��� _�������7� �    ?��� �����l��7� �    ?���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ��(~���׀        �  ��������        �  ��g�`����        �  �|_� <�����  �    ?�  ����<��;�  �    ?�  �S��|�_���  �    ?�  0����|�x�7�  �    �  ����� 8���  8�    �  �z�H�6���s��  <@    �  �������s�  .     �  �ސ�|���g��       ?�  ?�6�~������        ?�  ��������	��        �  {����և����        �  s����ȏ����        �  7���������  �    ��  ��������  �   ��� ����?���  ?�       ��� ������������ ���  ��� ��� ~����=�  �    ��� ���@~��  �       ��� �����>�����        �  �����>�����        �  ���4��������       �  ����������       �  ���������       ?�  #���������  �    �  ���?�����        �  9�?��??���  ?     ��  �~������  �   ��� ����?�����?�  ��   ��� ��1 ����?�  �    ��� ���?3����?�  �    ��� ������� � �    ��� ������    �       ��� ������@���� ���  ��� _�������/� �    ��� �����l��/� �    ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��~�`����            �|>� <�?���       �   �����<��;�  �    �   ��?�|�]|?�  \    ��  0����|�y�7� �   ��  ��������� ��   ��  �{���6���{�� �x   ��  �s�<������� �   ��  �w?��|������ ?�   ��  ?d�~����� �   ��� �������� �   ��� {���?և���?� ��   ?��� s���?ȏ���?� ��   ?��� 7����Ͽ���� ��  ��� ����������� =��  ��� �?�����~���� >��  ���� �]�����O��� M�  ���� �p7�~�C�� @�  ���� ��O� ~��?�?� �   ��� �ȟ�`>���� �   ?��� ��~~>�����  ~   ��� ���������� ��   ��� ������������ ���  ��� �y�����  �       ��� #���?��s��?� ��   ��� ���?��x  �       ��� 9� 9��>���       ��  �~���������  �    ��  ����������� �    ��  ��� ������ �    ��  ���s����� �    ��� ��?��� ?� �    ��� ������    ?�       ��� ������@���� ���  ��� _��?�����_� �    ��� ���?��l��_� �    ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��0`�0�       �� �}7� <���� �   �� ���D<��;� �   �� �7�l|�]��� �   �� 0��H|�y��7� �   ��� ������w� �   ��� �y�r6����}� �   ��� �}������| �   ��� �}�||����� �   ��� ?}�~����� �   ��� ������  �       ��� {�?��և� ��        ��  s����ȏ����        ?�  7����������        �  ����������  �    ��  ��  ��������       ��  ����B�����}� ��   ��� ����~��  ��       ��  �����~�����        �  �����>�����        �  ����>������       �  ������������  �    �  ����������  �    �  ����������  �    ?�  #���������  �    ?�  ���?�����        ?�  9߿��?����  ?     �  ���������  �    ��  ������������  ��   ��  ��� ������  �    ��  ���>�������  �    ��  ������ � �    ��� �����    �       ��� ������@���� ���  ��� _�������� �    ��� �����l��� �    ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��~�`����            �|~� <�����            ����<��;�            �x�|�_���            0����|�x�7�            ����� ���            �z�8�6������            ��8�������            ���|���g��        �  ?���~������  �    �  �����������  �    �  {����և�����  �    �  s����ȏ�����  �    �  7�����������  �    �  ��� ��������       �  ��� ��������        �  ���>��������        �  �����~���?��        �  �����~�����        ?�  �����>������  ?�    �  ��Á�>�����        ?�  ���������?��        �  �����������  �    �  ���������       �  #��������  �    �  ���?�����        ?�  9߿��?����  ?     �  ���������  �    ��  ������������  ��   ��  ��� ������  �    ��  ���?s����� �    ��� ������ � �    ��� �����    �       ��� ������@���� ���  ��� _�������?� �    ��� �����l��?� �    ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���o�����       �  ��K����?�F        �  ?| >������       �  |�
���i�        �  ~<�&���pi�        �  ��L>����qo�        �  ���5H8��?��        �  }�� (���� �^  `   ��  �  (~��  W�       ��� �  ���  w�       ��� ��  `�  ��       ��  �|  <� ��       ��  �� �< ;�        ��  � �|�_��        �  0���|�x 7�        �  � ��  ��        ��  �z| �6��| ��  c�   ��  �|  ���  |       ��� �y� <|��� ?� ��   ��� ?|  ~��  �       ��� �������	��        �  {�� �և����        �  s�� �ȏ����        �  7�� �������        �  ��� �������        ?�  ��� �������        ?�  ����������        ?�  ����~�����        ?�  ����~�����        �  ����>�����        �  ����>�����        �  ��� �������        �  ��<���<��  #�    ��  �~x ���x ��  t   ��  #�� ��|� �  �   ��� �� ?��|� � H �  ��� 9�` ��<` � � �  ��� �|  ���  �    �  ��� ��  ?���  ?�    @  ��� �   1 ��  ?�    @  ��� ��  ��   �       ��� �� ��� � �  ��� ��  �    �      ��� ��  �@   �      ��� _�  ��   �      ��� ��  �l   �      ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N>����qo�       �  ���5H8��?��        �  }�� (���� �^ �f   ��  �  (~��  W� �  ��� �  ���  w�       ��� ��  `�  ��       ��  �|  <� ��       ��  �� �< ;�        ��  � �|�_��        �  0���|�x 7�        �  � ��  ��        ��  �z| �6��| ��  c�   ��  �|  ���  |       ��� �y� <|��� ?� ��   ��� ?|  ~��  �       ��� �������	��        �  {�� �և����        �  s�� �ȏ����        �  7�� �������        �  ��� �������        ?�  ��� �������        ?�  ����������        ?�  ����~�����        ?�  ����~�����        �  ����>�����        �  ����>�����        �  ��� �������        �  ��<���<��  #�    ��  �~x ���x ��  t   ��  #�� ��|� �  �   ��� �� ?��|� � H �  ��� 9�` ��<` � � �  ��� �|  ���  �    �  ��� ��  ?���  ?�    @  ��� �   1 ��  ?�       ��� ��  ��   �       ��� �� ��� � �p  ��� ��  �    �      ��� ��  �@   �      ��� _�  ��   �      ��� ��  �l   �      ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ��(~���׀  �    �  �<������        �  ��x`��?��       �  �|s <����  
�    �  ���<�;�  �    �  �p�|�_��  �    �  0���|�x7�       ;�  ���� ��       =�  �z� �6�����       >�  �� �������       ?x  �� �|�����   �    ?�  ?��~�����        �  �������	��        �  {�� �և����        �  s�� �ȏ��?��        �  7�� �������        �  �� ������  �    ��  ��  ����  ��       ��  ��x B���x }�  g�  ��� ��  �~��  ��       ��  ����~�����        �  ����>�����        �  ����>�����        �  ����������        �  ���������        �  ��������        ?�  #�������        ?�  ��?�����        ?�  9ߜ��?���  �    �  �0 ����0��  (    ��  ��p ����p ��  |    ��  �x � ��x ��  $   ��  ��  ���  ��  x   ��  �  ��   �    �  ��� ��  �    �    �  ��� ��� �@� �     ��� _�  ��   �       ��� ��  �l   �       ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��~�`����            �|~� <�����            ����<��;�        `   �@�|�_A��  @     �   0�@�|�x@?7�  0     ��  ���� ���      ��  �z  �6�� ��  �@   ��  �|  ���� �     ��  �|  �|�� ��  `    ��  ?y  �~��  ��  �   ��  ��� ��� �       ��� {�  և�  �     ��� s�  ȏ�  �     ��� 7�  ?���  ?�      ��� ��  ?���  ?�     ��� ��  ?���  ?�  �   ?��� ��  ���  =� 	h   ?��� ��@ ~��@ =� �    ?��� ��� @~��� �      ?�� ��  `>��  � @   ��� ��� �>��� ��      ��  ��  ���  �  �    ��� ��� ?���� ?� x �  ��� �~  ���  �      ��� #�� ��|� �  ��   ��� �  ?��~  ��       ��  9ߜ��?���  �    �  �8 ����8��  4    ��  ��x ����x ��  d   ��  �p � ��p ��     ��  ��  ���  ��  x   ��  �  ��   �    �  ��� ��  �    �    �  ��� ��� �@� �     ��� _�  ��   �       ��� ��  �l   �       ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��~�`����            �|�8 <��8��  ��   ��  ���8�<�8;�  �   ��  ��8�|�^�8�  �   ��  0�� �|�x� 7�  �>   ��  �� �� � ��  �   ��  �z� �6��� ��  �   ��  �~� ����� �  �   ��  �~� �|��� ��  �   ��  ?~� �~��� ��  �   ��  ��� ���� ��  �   ��  {�  �և� ��        ��  s�� �ȏ����        ?�  7�� �������        �  ��  ���� ��        ��  ��  ����  ��       ��  ��� B���� }� �   ��� ��  �~��  ��       ��  ����~�����        �  ����>�����        �  ����>�����        �  ����������        �  ���������        �  ��������        ?�  #�������        ?�  ��?�����        ?�  9ߞ��?���  �    �  �8 ����8��  $    ��  ��x ����x ��  v   ��  �x � ��x ��  &   ��  ��  ���  ��  x   ��  �  ��   �    �  ��� ��  �    �    �  ��� ��� �@� � ��   ��� _�  ��   �       ��� ��  �l   �       ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��~�`����            �|~� <�����            ����<��;�            �x�|�_���            0����|�x�7�            ����� ���            �z�8�6������            ��8�������            ����|������            ?��~���q��       �  �������9��       �  {�� �և����       �  s�� �ȏ����  �    �  7�� �������  �    �  ��� �������      �  ��� �������       �  ����������  `    �  ���~�~�����       �  ����~�����        ?�  ����>�����  1�    �  ����>�����        ?�  ���L�������        �  �������?��        �  ��?����?��        �  #�������        �  ��?�����        �  9����?���  	�    ?�  ���������      �  ��8����8��  >    ��  �8� ��8��      ��  �� ��� ��  <    ��  �  ���   ��      ��  ��  ��    ��      ��  ��� ?�@� ?� ��@  ��� _�  ?��   ?�    @  ��� ��  ?�l   ?�    @  ���                                                                                                                                                                                                                                                                                                                                                                                 / / ����x���� �            ���������            �������?�F            ?| >�������            |�
����i�            ~9�&����i�            ��N�����qo�            ���uH8�����            }���(������^            ���(~����׀            �<�������            ��~�`����            �|~� <�����            ����<��;�            �x�|�_���            0����|�x�7�            ����� ���            �z�8�6������            ��8�������            ����|������            ?���~������            �����������            {����և�����            s����ȏ�����            7�����������            ������������            ������������            �����������            �����~������            �����~������            �����>������            �����>������            ������������            �����������            ����������            #��������            ��o?������            9�����?����            ����������            �����������            ���� �����            ��������?��            ��������            ������  `��            ������@  ��            _������  ��            ������l  ��                                                                                                                                                                                                                                                                                                                                                                                            / / ���� � ~���������      ���  ?���������      ���?�F �?���������      �����������~������      ����i�������������      ����i���Ǐ��������      ��qo�� ���N������      ������ ���������      �����^�  ��������      ����׀�Y ��������      �������c���~������      ����� ����������      ������Á@��������      ��;��� ��������      �_���������������      �x�7���� ��������      � ������p�2������      ������ �?��������      ����� �8��������      ������ � �������      ��������  �������      ������  ? ~������      �������  ? >������      �������   6������      �������   ������      ������p  ?  ������      ������   ?  ������      �����   �? ������      ������   ?�������      ������    ?�������      ������   �������      ������   ~�������      ������   3  ������      ������    � ������      �������  � ������      ���������������      ������� �� ������      �?������ r� ������      ��������  ������      ����� � ������      ��������������      ��?��?��������      �������� ������        `������  ������      @  ������  ������      �  ������  ������      l  ������  ������                                                                                                                                                                                                                                                                                                                                                                                      