�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                               ��                               ��                               ��                               ��                               ��                               ��                               ��              ����������������@��    `  0                    ���    `  0                    ���    `  0                    ���    `  0                    @��  0    0                    s���  0    0                    s���  0    0                    s���  0    0   ����������������@��  0    0                    y���  0    0                    y���  0    0                    y���  0    0                    @��Ǚ�>o�Ͱ                    |���Ǚ�>o�Ͱ                    |���Ǚ�>o�Ͱ                    |���Ǚ�>o�Ͱ   ����������������@�flٰ3;m�m�                    ~>�flٰ3;m�m�                    ~>�flٰ3;m�m�                    ~>�flٰ3;m�m�                    @�flٰ33m��0                    ~>�flٰ33m��0                    ~>�flٰ33m��0                    ~>�flٰ33m��0   ����������������@��lٰ?3m�g0                    |���lٰ?3m�g0                    |���lٰ?3m�g0                    |���lٰ?3m�g0                    @�6l۰a�m�m�                    y��6l۰a�m�m�                    y��6l۰a�m�m�                    y��6l۰a�m�m�   ����������������@�7Ǐ�a�m��                    s��7Ǐ�a�m��                    s��7Ǐ�a�m��                    s��7Ǐ�a�m��                    @�                               ��                               ��                               ��              ����������������@�                               ��                               ��                               ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �����?���������������������������������?���������������������������������?�����������������������������   �  `�                       ���������g����������������������������������g����������������������������������g��������������������������      a�x                       ����������������������������������������������������������������������������������������������������������  <    `                       ���Ã 8d������������������������������Ã 8d������������������������������Ã 8d����������������������������  <|�Ǜ`                       �����$�$�����������c��3����������������$�$�����������c��3����������������$�$�����������c��3������������  fv�`�`0                       �����$�1������������u�������������������$�1������������u�������������������$�1������������u���������������  ff�g�``                       �����$�1�?����������V����������������$�1�?����������V����������������$�1�?����������V������������  ~f�l�`�                       ���<�$�$�����������}U����������������<�$�$�����������}U����������������<�$�$�����������}U��������������  �f�l��                       ���<�$�$�����������v�����������������<�$�$�����������v�����������������<�$�$�����������v���������������  �f�g�a�                       �������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ������������������������������W���������������������������������W���������������������������������W����                                 �������������������������������������������������������������������������������������������������������                                 ���{���������������������������������{���������������������������������{�������������������������������                                 ���{����������������4��t�8�}�T������{����������������4��t�8�}�T������{����������������4��t�8�}�T����                                 ���zc��'͡�����������W[��V�Z��U������zc��'͡�����������W[��V�Z��U������zc��'͡�����������W[��V�Z��U����                                 ����u��ݮ����������W�{�V�Z��U�������u��ݮ����������W�{�V�Z��U�������u��ݮ����������W�{�V�Z��U����                                 ���~�u��ݮ���������u�W�x7V�Z��U������~�u��ݮ���������u�W�x7V�Z��U������~�u��ݮ���������u�W�x7V�Z��U����                                 ���~�u��ݮ���������u�WZ��V�Z��U������~�u��ݮ���������u�WZ��V�Z��U������~�u��ݮ���������u�WZ��V�Z��U����                                 ���~�u���n��������+�7X���V�k�V������~�u���n��������+�7X���V�k�V������~�u���n��������+�7X���V�k�V����                                 ���~���������������������������������~���������������������������������~�������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �������������������������������������������������������������������������������������������������������                                 �����������������?������8��q���������������������?������8��q���������������������?������8��q�����                                 ���{���������������������]w���������{���������������������]w���������{���������������������]w�������                                 ���{����������������������]w���������{����������������������]w���������{����������������������]w�������                                 ���zc��'���a��>��������]w���������zc��'���a��>��������]w���������zc��'���a��>��������]w�������                                 ����u����_������7]�멿�]w�ۮ��������u����_������7]�멿�]w�ۮ��������u����_������7]�멿�]w�ۮ�����                                 ���~�u����\.��~���]��뫿w]w����������~�u����\.��~���]��뫿w]w����������~�u����\.��~���]��뫿w]w��������                                 ���~�u����[�������]��뫾�]w�{��������~�u����[�������]��뫾�]w�{��������~�u����[�������]��뫾�]w�{������                                 ���~�u����[�������]��+��]w����������~�u����[�������]��+��]w����������~�u����[�������]��+��]w��������                                 ���~�����\!��>��8�������q�������~�����\!��>��8�������q�������~�����\!��>��8�������q�����                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������                                 ���������������������?��������������������������������?��������������������������������?������������                                 �������������������������������������������������������������������������������������������������                                 ���~4�v8c���������͏���������������~4�v8c���������͏���������������~4�v8c���������͏�������������                                 ����]w�]����������~�w����������������]w�]����������~�w����������������]w�]����������~�w�������������                                 ���~]vA��������������������������~]vA��������������������������~]vA������������������������                                 ���}�]u�_���������������������������}�]u�_���������������������������}�]u�_�������������������������                                 ���}�]e�]���������ˮ�w���������������}�]e�]���������ˮ�w���������������}�]e�]���������ˮ�w�������������                                 ���a�c��������p͏���������������a�c��������p͏���������������a�c��������p͏�������������                                 �������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �����������������8a�>����������������������������8a�>����������������������������8a�>������������                                 �����������������׮��������������������������������׮��������������������������������׮����������������                                 �����������������׮��������������������������������׮��������������������������������׮����������������                                 ���|N5�����������׮���;DÌ���������|N5�����������׮���;DÌ���������|N5�����������׮���;DÌ�������                                 �����������������7����[]�������������������������7����[]�������������������������7����[]���������                                 ���}�������������׮����{[]����������}�������������׮����{[]����������}�������������׮����{[]��������                                 ���}��������������׮���#�[]u����������}��������������׮���#�[]u����������}��������������׮���#�[]u��������                                 ���}��������������׮������]u����������}��������������׮������]u����������}��������������׮������]u��������                                 ���������������8a�Y�=�C����������������������8a�Y�=�C����������������������8a�Y�=�C��������                                 �������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        