�P  �G� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  �                        ����� ��                        ����� ��                        ����� ��                               ��                        ����� ��                        ����� ��                        ����� ��              ��������� ���@� 0                  ����� �� 0                  ����� �� 0                  ����� �� 0                  �    @�       0            ����� s��       0            ����� s��       0            ����� s��       0  ������������@�       0            ����� y��       0            ����� y��       0            ����� y��       0            � �  @�7�������;<��         ����� |��7�������;<��         ����� |��7�������;<��         ����� |��7�������;<���������������@����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         ����� ~>����6��l�ٳf�         � �� @���������3f��         ����� ~>���������3f��         ����� ~>���������3f��         ����� ~>���������3f���������������@����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         ����� |�����3�����3f�`         � �  @�0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͰ         ����� y��0ٶ�6��l�ٳfͿ������������@�0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         ����� s��0ٶ�������<��         �    @�                        ����� ��                        ����� ��                        ����� ��              ��������� ���@�                        ����� ��                        ����� ��                        ����� ��                               @�                                 �                                 �                                 �              ������������������                                 �                                 �                                 �                                 �                                 �                                 �                                 �              ����������������  ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ��                               ���                               ���                               ��?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������8�1�������[S�Ɵg�f�������������8�1�������[S�Ɵg�f�������������8�1�������[S�Ɵg�f����������?�������������������������������������{~���u��w���Mw�o[�Z�������������{~���u��w���Mw�o[�Z�������������{~���u��w���Mw�o[�Z���������?�������������������������������������{p���u����]w��o�n��������������{p���u����]w��o�n��������������{p���u����]w��o�n����������?��������������������������������������n���u�����]w��w�v��������������n���u�����]w��w�v��������������n���u�����]w��w�v���������?�������������������������������������{n���u��wݺ�]w��[�Z��n������������{n���u��wݺ�]w��[�Z��n������������{n���u��wݺ�]w��[�Z��n��������?��������������������������������������p����_����]���g�f��������������p����_����]���g�f��������������p����_����]���g�f���������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������o�������o������������������������o�������o������������������������o�������o����������������������?�����������������������������������o�������o�������������������������o�������o�������������������������o�������o�����������������������?�����������������������������������)�ʉ�c1�)����S��3i���-���������)�ʉ�c1�)����S��3i���-���������)�ʉ�c1�)����S��3i���-�������?�����������������������������������f�ڶ�}n��f��[��w������k����������f�ڶ�}n��f��[��w������k����������f�ڶ�}n��f��[��w������k��������?�����������������������������������n�ڶ�a`��n��[����.�U�g����������n�ڶ�a`��n��[����.�U�g����������n�ڶ�a`��n��[����.�U�g��������?�����������������������������������n�ڶ�]o��n����������U�k���������n�ڶ�]o��n����������U�k���������n�ڶ�]o��n����������U�k�������?�����������������������������������n�ڶ�]n��n��[��w������m����������n�ڶ�]n��n��[��w������m����������n�ڶ�]n��n��[��w������m��������?�������������������������������������ڶ�a�������]��7n���n�����������ڶ�a�������]��7n���n�����������ڶ�a�������]��7n���n�������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������?������������������������������������4��|�c0��3��}�2ߌ��N?��������4��|�c0��3��}�2ߌ��N?��������4��|�c0��3��}�2ߌ��N?�����?�����������������������������������u�]齚�}n��t���u�齵ֿ����5��������u�]齚�}n��t���u�齵ֿ����5��������u�]齚�}n��t���u�齵ֿ����5������?�����������������������������������u�A뽺an����}��U����t�������u�A뽺an����}��U����t�������u�A뽺an����}��U����t�����?�����������������������������������u�_뽺�]n��}���}���Uֿu���u��������u�_뽺�]n��}���}���Uֿu���u��������u�_뽺�]n��}���}���Uֿu���u������?�����������������������������������u�]뽺�]n��u���u�����u���u��������u�]뽺�]n��u���u�����u���u��������u�]뽺�]n��u���u�����u���u������?������������������������������������7c뾻ap�������6���v?��������7c뾻ap�������6���v?��������7c뾻ap�������6���v?�����?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������������������}���������������������������������}���������������������������������}�������������������?�����������������������������������������������}���������������������������������}���������������������������������}�������������������?�����������������������������������c�9��1�|�1��<�϶�[���m����������c�9��1�|�1��<�϶�[���m����������c�9��1�|�1��<�϶�[���m��������?�����������������������������������]t��]n����n��}�������}�������������]t��]n����n��}�������}�������������]t��]n����n��}�������}�����������?�����������������������������������_u��_n���n��}�ߪ���a𫪿���������_u��_n���n��}�ߪ���a𫪿���������_u��_n���n��}�ߪ���a𫪿�������?�����������������������������������_u��_n�}��n��}�諸�������������_u��_n�}��n��}�諸�������������_u��_n�}��n��}�諸�����������?�����������������������������������]u��]n����n��}��ݺ��]���������]u��]n����n��}��ݺ��]���������]u��]n����n��}��ݺ��]�������?�����������������������������������c���cq�~����~��������w���������c���cq�~����~��������w���������c���cq�~����~��������w�������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������7y��68Ϗ�c6��vq�_	��Nc�����������7y��68Ϗ�c6��vq�_	��Nc�����������7y��68Ϗ�c6��vq�_	��Nc��������?�������������������������������������{w���_���]v�_u��^���5��uo����������{w���_���]v�_u��^���5��uo����������{w���_���]v�_u��^���5��uo������?�������������������������������������{w�߇�Av�_v�^�Uu��u�����������{w�߇�Av�_v�^�Uu��u�����������{w�߇�Av�_v�^�Uu��u�������?�������������������������������������{w����w��_v�_wo�^�uUu��u�����������{w����w��_v�_wo�^�uUu��u�����������{w����w��_v�_wo�^�uUu��u�������?�������������������������������������{w���_w��]y�_e��^�v�u��uo����������{w���_w��]y�_e��^�v�u��uo����������{w���_w��]y�_e��^�v�u��uo������?������������������������������������9}��68��c��ߖq�_��vc�����������9}��68��c��ߖq�_��vc�����������9}��68��c��ߖq�_��vc��������?������������������������������������������������������������������������������������������������������������������������������������������?�����������������������������������?����������������������?�����������?����������������������?�����������?����������������������?���������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������}��������������������������������}��������������������������������}�����������������������������?���������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������?�����������������������������������mMc�8�u?i�?|�cm��2|ko���������mMc�8�u?i�?|�cm��2|ko���������mMc�8�u?i�?|�cm��2|ko�������?�����������������������������������m5]��{t�릶��齚�]mu�����o���������m5]��{t�릶��齚�]mu�����o���������m5]��{t�릶��齚�]mu�����o�������?�����������������������������������UuA��{u�����~뽺]U��*����������UuA��{u�����~뽺]U��*����������UuA��{u�����~뽺]U��*��������?�����������������������������������Uu_���u�����뽺�]U}��������������Uu_���u�����뽺�]U}��������������Uu_���u�����뽺�]U}������������?������������������������������������u]��{e�뮶��뽺�]�u����������������u]��{e�뮶��뽺�]�u����������������u]��{e�뮶��뽺�]�u�������������?������������������������������������uc�����n�?��c���7|+�����������uc�����n�?��c���7|+�����������uc�����n�?��c���7|+��������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������������������������������������������������������������������������������������������������������?������������������������������������47X�~3�q�c�~3f8���������������47X�~3�q�c�~3f8���������������47X�~3�q�c�~3f8������������?�����������������������������������m���_Z��ٮ��mu������������������m���_Z��ٮ��mu������������������m���_Z��ٮ��mu����������������?�����������������������������������m���XZ��۠��m��,��������������m���XZ��۠��m��,��������������m���XZ��۠��m��,������������?�����������������������������������mu��WZ��ۯ��m}������������������mu��WZ��ۯ��m}������������������mu��WZ��ۯ��m}����������������?�����������������������������������mu��WZ��ۮ��mu������������������mu��WZ��ۮ��mu������������������mu��WZ��ۮ��mu����������������?�����������������������������������m��9Xk�7���m�~768_��������������m��9Xk�7���m�~768_��������������m��9Xk�7���m�~768_������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                ����������������������������������������������������������������������������������������������������������?������������������������������������������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                 ����������������������������������������������������������������������������������������������������������                                                                                                                                          �����������������������������������                                                        