�P   ˀ� �Ƿ���?�����?������������������?�����?����������������x                        D������� �� _������   ������ �� _������   �H                           >     �������     ?������     �������     ?�������                           8N     �     �     8          �     �     8     �                        �{������?������� /�����������?������� /��������                        B9��������_������� w���������_������� w��                            >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     D                        ���������������{�~/�����������������{�~/�������                        �9�������^�������? `u�������^�������? `t�                            >     �������     ?������     �������     ?�������                           @N     �     �     8          �     �     8                             �|���}��� �?��������, ������}��� �?��������, ������                        P� ��������P >������ 5 ��������P >������ 4�                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     4                        ��7��?y��� 0?��������� �����?y��� 0?��������� �����                        H8  ������� @ ������   ������� @ ������ �                           >     �������     ?������     �������     ?�������                            �     �     �     8          �     �     8                             ��������  ?���������  ��������  ?���������  �����                        Q8�  ������  H  ������  �  ������  H  ������  �                           >     �������     ?������     �������     ?�������                            N     �     �     8          �     �     8                              ���������  ?���������  ���������  ?���������  �����                         9�  ���_���  \  ������  �  ���_���  \  ������  �                            >     �������     ?������     �������     ?�������                           N     �     �     8          �     �     8                              �{�'��i���  ?��������` ���'��i���  ?��������` �����                        8�  ������ M� ������X �  ������ M� ������X ��                           >     �������     ?������     �������     ?�������                           �N     �     �     8          �     �     8     D                        �������������������������������������������������������                        8           @                     @          �                           ?���������������������������������������������������                           O�������������������������������������������������� $                        �o�                                                 ��                        ;����������������������������������������������������                           ?���������������������������������������������������                           �O��������������������������������������������������	                        ������������������������������������������������������x                         8           @                     @          �                            ?���������������������������������������������������                           O�������������������������������������������������� �                        �������������������������������������������x                        �8 ���}����cA��������4 ���}����cA��������4�                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8     �                        ������>���w�|��������������>���w�|�������������                         8  ��������@ �������84  ��������@ �������84�                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ������ ����e����������[����� ����e����������[����                        8 ��}����#@��������4 ��}����#@��������4�                            ?�������     �������     �������     �������     �                           @N     �     �     8          �     �     8                             ������������\�����8��������������\�����8������x                        9���������X��������5���������X��������4�                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      �                        ��������ꏾ������>���8|�[�����ꏾ������>���8|�Z��                        9�������x4�\������O��������x4�\������O��@                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                              ���������������?(�����;������������?(�����:��                        %9������x4�\8��������O�������x4�\8��������O��P                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �?���~��~���_H�����-����u���~��~���_H�����-����u���                         9����?�߸��\ 9�������}�����?�߸��\ 9�������}��                            ?�������     �������     �������     �������     �                           �N     �     �     8          �     �     8                             ���/���o������������O���A�/���o������������O���A���                         9��������_�`_�п����5��������_�`_�п����4�                            ?�������     �������     �������     �������     �                           RN     �     �     8          �     �     8     $                        �Ϸ����������P����������E����������P����������E
��                         9� ��A����_� ��������� ��A����_� ���������                            ?�������     �������     �������     �������     �                           0N     �     �     8          �     �     8                             ����������S�?�����(��7�C��������S�?�����(��7�C���                        b�����q�����_�+ ����������q�����_�+ �������(                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      T                        �����������~������h��y�G���������~������h��y�G���                         9�����s����_�~8��?���������s����_�~8��?�����                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ������?���O��?����/���� z���?���O��?����/���� z��                        �9���� �����_�<����������� �����_�<��������                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      d                        �߶������?_������������������?_��������������                        �9�����_����_�p(�Pu����������_����_�p(�Pu������@                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                             ��?��w���@�������$�!�?��w���@�������$�!���                         ����������_o��Pp��������������_o��Pp������                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                             ��̿�'���<?�>���������c�̿�'���<?�>���������c��x                        �����s/����_����W2�?�������s/����_����W2�?����(                           ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8     �                        ������o��C�o�>�� ����?��C����o��C�o�>�� ����?��C���                        P9���A�w����[����W{�?������A�w����[����W{�?����                            ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              ���� ������_�f�� ��������Fk� ������_�f�� ��������Fj��                         9�����e����\_���W� >�������e����\_���W� >���                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8      4                        ����������`y���������Ǒ���������`y���������Ǒ���                         8
�������@�������?�t
�������@�������?�t�                            ?�������     �������     �������     �������     �                           N     �     �     8          �     �     8                             ���������������������9���������������������9�����                        �� q������@�����?�4 q������@�����?�4��                           ?�������     �������     �������     �������     �                            N     �     �     8          �     �     8                              �߷��������~>������o��������������~>������o��������                        �8  ����3��@ �����?�  ����3��@ �����?���                           ?�������     �������     �������     �������     �                            N    � �  �  p  8        � �  �  p  8                            ������c���������v?�)���w�����c���������v?�)���w����                        9� ~������X w����ݏ�� ~������X w����ݏ��                            ?������ �  ���w���    ������ �  ���w���    �                           N  � � �  �  �  8  >    � � �  �  �  8  >   D                        �6������������?����7��������������?����7����                        9� � ������_� ���?����e� � ������_� ���?����d�                           ?������ �  �������  >  ������ �  �������  >  �                           ��  � � �  � �  8      � � �  � �  8                            ���ߟ�ҽ���������+��~���ߟ�ҽ���������+��~����                        9� � }C�����_����?��E� � }C�����_����?��D�                           ?��ߟ��� �  �������  ~  ��ߟ��� �  �������  ~  �                           �N  ?� � �  � �  8  ��   ?� � �  � �  8  ��                         ����ߟ��������������~�K�ߟ��������������~�J��                        9� � mG�����_�������� � mG�����_��������                            ?��ߟ��� �  �������  ~  ��ߟ��� �  �������  ~  �                           AN  ?� � �  � �  8  ��   ?� � �  � �  8  ��                         �����ߟ���������������~���ߟ���������������~����                         9� � g�����_ �� V���� � g�����_ �� V����                            ?��ߟ��� �  �������  ~  ��ߟ��� �  �������  ~  �                           N  ?� � �  � �  8  ��   ?� � �  � �  8  ��  4                        ���������� ���������0���������� ���������0����                        8� � �����N �� ����� � �����N �� �����                           ?������    �������  0  ������    �������  0  �                           �N  ?� � �  � �  8  ��   ?� � �  � �  8  ��                         ������?����� ���������������?����� �������������x                        8  � �����@  �� ������  � �����@  �� �������@                           ?���?���     ������     ���?���     ������     �                           N  � � �  � �  8      � � �  � �  8     �                        �����������a�������������������a�������������                        F8  ~�����@  p'�������  ~�����@  p'��������`                           ?������     ������     ������     ������     �                            N  � � �  �  �  8  >    � � �  �  �  8  >                           ��7���������a?���w�����������������a?���w����������                        �8   ����@   '�������   ����@   '��������                            ?������     ������     ������     ������     �                            �  � � �  �  �  8  >    � � �  �  �  8  >                           �}������������?�����������������������?��������������                        !8    ����@   ��� ?��    ����@   ��� ?���                           ?������     ��� ���     ������     ��� ���     �                           �N  � � �  � �  8 ��   � � �  � �  8 �� $                        �߷���������p��������������������p�������������                        8  �?������@ �#�������  �?������@ �#��������`                           ?������ �  ������ �� ������ �  ������ �� �                            N  �� � ?�  � �� 8 ��   �� � ?�  � �� 8 ��                         �߷�������������p��������������������p���������                        8   �����@   �8�� ?��   �����@   �8�� ?���`                           ?������     ��� ���     ������     ��� ���     �                            N  � � �  � �  8 ��   � � �  � �  8 ��                         ����������������w������g���������������w������g����                        8@  f ����D  ` ������@  f ����D  ` �������                           ?������     ������     ������     ������     �                            N  � � �  �  �  8  >    � � �  �  �  8  >                           ��7��������Ͽ����w�����������������Ͽ����w�����������                         8  A �����@  t ������  A �����@  t �������                            ?������ �  ���w���    ������ �  ���w���    �                           "�  � � �  �  �  8  >    � � �  �  �  8  >  ,                        ������?���?��������������������?���?�������������������                        �� � �����@p � ������ � �����@p � �������                           ?���?��� �  �������  8  ���?��� �  �������  8  �                           N  � � �  � �  8      � � �  � �  8     $                        �����������ǿ���������|{����������ǿ���������|{����                        �9��� ~?����[�� �������� ~?����[�� ������                            ?������ �  �������  |  ������ �  �������  |  �                           @N  ?� � �  � �  8  ��   ?� � �  � �  8  ��                         ����������������������9���������������������9���x                        49�� �~?���]�   �� ?���� �~?���]�   �� ?���@                           ?������     ��� ���     ������     ��� ���     �                           N  � � �  � �  8 ��   � � �  � �  8 ��  �                        ���~7����ߌ���������������~7����ߌ����������������                        
9��� ����X��P �������� ����X��P ������                           ?��~��� �  ������ �  ��~��� �  ������ �  �                           N  �� � ?�  � �� 8 ��   �� � ?�  � �� 8 ��                         ���������?������������g��������?������������g����                         8 �� �����@p�  ������ �� �����@p�  �������                            ?������ ?�  ����?�� �  ������ ?�  ����?�� �  �                            N �� � �  � �� 8 ��  �� � �  � �� 8 ��                          ���������������������w��������������������w����                        8�� ���@ �  W�������� ���@ �  W��������                           ?������ �  ������ �  ������ �  ������ �  �                           @N �� � ��� � ?�� 8 ��  �� � ��� � ?�� 8 ��                         �����������x���������7�w���������x���������7�w�
��                        8������@���������������@����������P                           ?������ �  ������ �  ������ �  ������ �  �                            N �� � ��� � ?�� 8 ��  �� � ��� � ?�� 8 ��                          �7��~��������������������~��������������������                        8���x��?�G����׀o������x��?�G����׀o����`                           ?��� ��� �   ������ �  ��� ��� �   ������ �  �                           �� �� ���� � �� 8 ��  �� ���� � �� 8 ��                         ��� ����������� 8?�������� ����������� 8?����������                        "9���  @ � ?�_���  � ������  @ � ?�_���  � ����                            ?��� ��� �   ��� ��    ��� ��� �   ��� ��    �                            N �� ���� � �� 8 ��  �� ���� � �� 8 ��                          ��� ����������� ?���������� ����������� ?�����������h                         9��       ?�_�       ����       ?�_�       ���                            ?��  ���     ��  ��     ��  ���     ��  ��     �                           	N �� ���� � ��� 8 ?��  �� ���� � ��� 8 ?��  �                        �������������� ��������������������� ������������                        (9����  ����_���  ��������  ����_���  �����                           ?��������� ������ �� ��������� ������ �� �                            N ������� � ��� 8 ?��  ������� � ��� 8 ?��                          ����?������� �����������?������� �����������                        9��� p���W��   ������ p���W��   �����                           ?��� ���   �� �� �  ��� ���   �� �� �  �                           N ������� � ��� 8 ?��  ������� � ��� 8 ?�� $                        �6��?������������������?������������������                        9���� 6���_��  `������� 6���_��  `����                           ?��� ���   �� �� �  ��� ���   �� �� �  �                           �� ������� � ��� 8 ?��  ������� � ��� 8 ?��                         �������������������������������������������������������                        �           @                     @          �                           ?���������������������������������������������������                           O�������������������������������������������������� $                        ���                                                 ��                        �����������������������������������������������������H                           ?���������������������������������������������������                            O��������������������������������������������������                         �������������������������������������������������������                        �8           @                     @          �                            ?���������������������������������������������������                            O��������������������������������������������������                         ������������c��!��/����;�� �������c��!��/����:��                         ������ ?x�_�����`�������>� ?x�_�����`�����                           >     �������     ?������     �������     ?�������                            N     �     �     8       � �     �     8                              �����������������]�/����8;��������������]�/����8:��                         9���>  ��_������ �������>  ��_������ �����                            >     �������     ?������    �������     ?�������                           �N     �     �     8       � �     �     8                             �ݷ�����������#���Yo�/����;����������#���Yo�/����:��                        	9��� � @��_������������ � @��_����������                           >     �������     ?������    �������     ?�������                           "N     �     �     8       � �     �     8     $                        ���~� }r������`�/����:~��}r������`�/����:��                        �9������`A����_����8��������σ�`A����_����8������                            >     �������     ?������  � �������     ?�������                            N     �     �     8       � �     �     8                              �o�>�,���x4������o���O�>��,���x4������o���O���                        9������pA����_���>�����������pA����_���>�������                           >     �������     ?������  � �������     ?�������                           �N     �     �     8       � �     �     8     	                        ���>�r�,N���x4����/������O�>�,N���x4����/�������O���                        A9������p@����_���? ����� ��p@����_���?<���                           >     �������     ?������    �������     ?�������                           N     �     �     8      � �     �     8      D                        ���?��}#��߸�߳����>+����}�?��=#��߸�߳����>+����}���                         ���~��}p x��'O���-�� ��t��g"�}p x��'O���-�� ��t�                           >     �������     ?������    �������     ?�������                           N     �     �     8      � �     �     8      $                        �������r������?��(��0�;�� �r������?��(�����:��                        8/���o��E�B�������>��/��o��E�B�������W���@                           >     �������     ?��0��    �������     ?�������                           N     �     �     8 ��  �� �     �     8      $                        �������QB����믯���,���������QB����믯���,�������                        9�����  �P�������������.�  �P������  ���                            >     �������     ?������ �� �������     ?�������                           DN     �     �     8 ��  ����     �     8     D                        ��;�M�P���������ԏ���k\�
;�/�����?������������
��                        �9����� ���\������������/ � �\�����
����                            >     �������     ?��c��     ���?���     ?�������                           N     �     �  p  8 ?��  ���� �  �     8     D                        �߶38x�������3�s��?˿�32/���������3���?������                        ������1����\����W��������o1���\�����W�����X                           >     �������     ?�Ü���     ������     ?�������                            N     �     � �  8 ?��  ���� �  �     8                             �����`0��������������_�������������������������                         8�`0?��@��@?���������?��@ �@?�����  ���                            >     �������     ?�� ��     ������     ?������                            N �� �     � �  8 ��  �� � �  �     8 <                          �����o� z�_����/����u�_������ z�_�����/����u������                         8{o2��� ��A��x������x�������A�������<��                            >   ������  x  ?�� ��     �������     ?������                           N �� � �   � �  8 ��  �� � �  � 8   8 <                          �=�����z�`����������p�/����ȋ�z����������p������                         8;o2w�}�`��A��������'�<tw�}����A��?���ͼ��                            >   ��`����  �  ?�� ��     �������    ?������                           �N �� � �   � �  8 ��  �� � �  � ?�  8 < $                        ���3Bo����.n���4
|}��2�/���3@�����/����4����2�>П��x                         9̻2'��� �\��~b����'�̼t'�����\˯�������                            >   ��.���  |  ?�� ��     ������� �  ?������                           N �� ���  � �� 8 ��  �� � �  � �  8 <  �                        ��6a
������Ǜ���<y�{����aE�����������{�>����                        9��o�o����]� >f�����G���:o�o����]�/������<��                           >   �������  <  ?�� ��     ������� #�  ?��<���                           0� �� ���  � �� 8 ��  �� � ?�  � �  8 ��                         ��;�������������a�����;������a����8�����3����                         ������q}���_�~�������� ����q�|�_�~���������                           > �  �������   ?������  �� ���a��� 8|  ?������                           N �� ���  � �� 8 ��  �� � ?�  � ��  8 ��                         �������n���}���W�F������{�����n���%���w�F����3�z��                         ������� A����_�����   ���  �� B�9��_����/����                           > �  ���=��� �  ?�� ��     ���!��� w�  ?������                           N �� ���  � �� 8 ��  �� � ?�  � ��� 8 ��                          ��7�������Ϟ������o�����;�������ׅ���s��o���3�:��                         9����� C���_������������x @9��_����������                            > �  ��ώ��� �  ?������ �� ������ s� ?������                           @� �� ���  � �� 8 ?��  ���� ?�  ���� 8 ��                         ����������������������������8����K������������3���                         9����� C���_�����P�������? @���_�����P����                            > �  ������ �  ?������ �� ������ ��� ?������                           N �� ���� � �  8 ��  ���� �  ���� 8 ��  T                        ���~������?�?������������
~���~���������������3�
��                        $9�����`F� _���?��������`@�_���������@                           > �  ��?�?��     ?������ �� ������ ��� ?������                            N �� ���� � �  8 ?��  ���� �  ���� 8 ��                          ����������?��ƿ����h?��k�������t�ƿ}����h?����j�x                         8�  �~��?@��a?��   ��  �~ ��?@���o��   ��                            >     ��?����     ?�� ��     ��������` ?�� ���                           N �� ���� � �  8 ��  �� � �  ���� 8 ��  �                        �������������������?�?�J�������������y����?����J��                        9� ��~���P�����  8�����~  �P���g��  ��                           >     �������     ?�� ?��     �������` ?�� ���                            N �� ���� � �  8 ��   � � �  ���� 8 ��                          �����������������x�,�?���������������z�>g�,�?���x                        9����~���Q������  8�����~  �Q�������  8��                           >     �������     ?�� ?��     �������>` ?�� ?���                           N  � ���� �  �  8 ��   � � �  ���� 8 ��  �                        ��6o������������������?��o�������������>w������p                         9�����|���Y������ |8 �����| � Y�������  x �                            >     �������  �  ?�� ?��     �������>0 ?�� ���                           �  ?� �?��� � �� 8 ��   � � �� ���� 8  �� �                        ����?�������������O���������0a����?�?�����w����������                        9��?���8��� _�����Ӏ � ��?���8 ?�  _����Ӏ �� �P                           >  ?� ������� �@ ?�����  0  ��?�?���>0 ?�������                            N �� �?��� � ?�� 8 ��   �� � ��� ���� 8 ��                          ����� ����������������������8a���������������� ����                         9������ ?q�� _�� ��  � ��?���      _��7�� �� �                            >     ��q����     ?�����  8  ��  ���~0 ?�� ���                            N �� ���� � �� 8 ��   �� ���� ���� 8 ��                          �������������������_��������<e������^���~�_���������                        P9������ '��߀_������  �	���?���  ��߀_���7�� ����                            > �� ������� ?� ?�����  <  ����_��	�~0 ?�������                           N �� ���� � �� 8 ��   �� ���� ���� 8 ��  D                        ���������������� O��������<%����������O���>����                         9�� �� !����_�����  �	���?���  ���_�a�7��   ��                            >     ������ �  ?�����  <  ����� �0 ?�� ���                           �N �� ���� � �� 8 ��   �� ���� ���� 8 ��                         ��7��￀���'���������������|3�����?���������������                        �9���?�� ���_�� �� �������    �_���g��   ��                            >     �����     ?�����  |  ��  ?����` ?�������                           �  � �?��� � ?�� 8 ��  �� � ��� ���� 8                             �������~��O�����������������|1�~���������l���������                        9���?�� ?���_�� ��� �������    ��_������   ��`                           >     ������     ?�����  |  �������` ?�������                            N  � ���� � �  8 ��  �� � �  ���� 8                             �������~��??�����?����������~3�~���������O����������                         9�����  � �_�� ��� � �����    �_�����  >��                            >    ��??��     ?�����  ~  ������ �@ ?�������                            N  � ���� � �  8 ��  �� � �  ���� 8                             ���������������������������������������?������������                        ������ ��� _������    �� �� � _�?����  >� �                           >    ������� �  ?�� ��     ������ ?�� ?�������                            N  � ���� � �  8 ��  �� � �  � ��� 8                             ������������������������'���������������������|����                         ������� ��� _������ �� ������  �@ _������  ? �                           >    ������� �  ?�����  �  ������ ��� ?��<���                           N  ?� ���� � �  8 ��  �� � �  ���� 8  ��                          ��7����������?�����o�����#��������������?������������                        �9�������    _������� ��������@ _�  �� ? �                            >  � ��  ?�� �  ?����� �  ������     ?��>?���                           �  � ���� � �� 8 ��  �� � �  � ��� 8 ��  ,                        ���G?�����9�����s��/�/���1��G3���?�����r���/��������                        �9������o����_���?����� 5�����o��@_������  4�                            >  � ������� �  ?����� �  ������� �� ?��~?���                           N  � ���� � �� 8 ?��  ���� ?�  ���� 8 ��  D                        ��'?����<��?��s��'�����9��'3���?�����s?�����������x                        �9�����w�    _�� ?���� �����w�  ` _�  ��   �                            >     ��  ?��     ?����� �  ��� ���     ?�� ?���                           N  � ���� � �� 8 ?��  ���� ?�  � ��� 8 �� �                        ���s�~2��� ���;������8��s��?������;�/����������                        9����c�?�@ _�����?�� �g��?�c��@ _���?��?� ��                           >  ~  ��  ��� �  ?��� �� �  ������     ?������                            N  �� � ��  � �� 8 ��  ���� �� � ?�� 8 ��                          ����������~������������x�����?���?�?���߃������o���x                        9��������� _������� ����?��?�  _���?���� �`                           >  �  ��~ ��� �  ?��� �� �  ��?�?�� �  ?������                           N �� � ��  � ?�� 8 ��  ���� ��� � ?�� 8 ��  �                        �������������ߟ�������������>?���ǟ��߿�������w����                        
������� ��� _������ ����?� �� _������� �                           > �  ������ �  ?��� �� �  ����� ?�  ?������                           N �� ���� � �� 8 ��  ������� � �� 8 ��                         ������~������� /�������~"�~�������� /���w���X                        �9���������_ߟ�����w�����?���_߿������w��                            > �  ��� �� �  ?��  �� �  ����� ?�  ?������                           N �� ���� � �� 8 ��  ������� � �� 8 �� �                        ��7���}����?������~/�0���� ���~�����~/�w������                        9��������^�����?�`u�� ����^������ `t�                           > �  ��� ?�� �  ?�0  �    ��~ ��    ?������                            � �� ���� � �� 8 ���� ?������� � ��� 8 ��                          ��6�������������8?��, ��?�������� ������p��, �����                        9 � ����  P ?����   5    O���  P ������  4�                            > �  ��� �� 8   ?�   ?�     ��� �� p   ?�� ���                           0� �� ���� � ��� 8���� ������� ���� 8 ��                         �������?��������?���� ������������ ����������� ������                         8    ?��    @   ������� ?�����    @   ����   �                            >     ��  ��     ?������ ?�����  ��     ?��  ���                           N ������� ���� 8���� ������� ���� 8 ��  t                        �������������������� ���?������������������ ?������                        8��������� H ����������?� o����� H��������� ��                           > ���������� ��� ?��� ?� ?�  ���������� ?�������                            N ������� ���� 8���� ������� ���� 8 ��                          �Z����?������������ ���?����������������� ?������                        9���?�_���  \ ���������?� o�_��� \�������  �                            > �  ��� �� �   ?��� ?� ?�  ��� ���   ?��� ���                           �N ������� ���� 8���� ������� ���� 8 �� 
T                        ��'��?�������~����`���?�'����������}����`?������                        8���?����  M����������?� o���� M��������  ��                           > �  ��� �� �   ?��� ?� ?�  ��� ���   ?��� ���                           N ������� ���� 8���� ������� ���� 8 ��                         �������������������������������������������������������                         8           @                     @          �                            ?���������������������������������������������������                           O��������������������������������������������������                         ��4                                                 ��                        ;����������������������������������������������������                           ?���������������������������������������������������                           !���������������������������������������������������                        �߰                                                  ��                         8                                                  �                            8                                                  �                            O��������������������������������������������������                        ���                                                  ��                         ?���������������������������������������������������                            ?���������������������������������������������������                           BO��������������������������������������������������$                        �������������������������������������������������������                        C?���������������������������������������������������0                           ?���������������������������������������������������                            @                                                                           ��?����������������������������������������������������                        ?���������������������������������������������������@                           ?���������������������������������������������������                            �                                                                           �������������������������������������������������������                         ?���������������������������������������������������                            ?���������������������������������������������������                           @                                                   $                        �������������������������������������������������������                        �����������������������������������������������������H                                                                                                                                                                                       ������}��������}�����ٻ���������������������������                           �   P@ ��  �@ H�   (P  � � ��   �                                                                                                            @�     �  &D "  �B  �   $ �@@ (�d                        ������������^�����}�����v�������������_o������������0                        �@��  ��@!�@` �      � � B   (	  � 	                                                                                                           �   �	   � $ (�  @�@B 	  ��         �                        �=��������߯}��߿��}�6����}���w���������������������                         @ �     D$de    �    PH A   D � @                                                                                                            @  P�  @��� �p " �  �@D @  	 A  ,                        ����������o�v�����������������y��������������a�����                          �     @A A �X��  ��!(  !@�  @�   �                                                                                                             � �S D� �   �          �@ h@ @ � �QB$                        �����������{~���������������?�W���������a�=����������x                        A�@   � @  "  � �   @ P�        �    �                                                                                                          @  @P	�� @%   ! "  �0�     � �hP@   P   �                        ����������~����������������_����ޗU���������|��������                          @��       @ @1PPH T       @ �  @@�                                                                                                          #    �     `  �  0	!h�   d$H �  !  T                        ������������������������������������������o�����~��                        � (  D d@ 
 K� H0   �P ���I   D	!@$ A  Ԅ BP                                                                                                          B0  (�   �   �!      �0   �  �                        ��}����������������_�?��������=����7�������g������x                        P1  �E@ h@ !      A  � � ` (@ �                                                                                                          H�  �       �� �B!  DC  �(�   @ �     �                        ��_߿���������������������_�?�������g�������������}�                          �B $	       B� 
 �  \�H �  *  H @                                                                                                            � @    H�! D     @� �     �         ��                        �                                                                                                                                                                                                                                              ������������������������������������������������������                        �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                             ������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            