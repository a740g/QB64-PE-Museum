�P  �>  P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �����                        �����    �����    �����    �����              �����    �����    �����              �����    �����    �����                        �����    �����              �����    �����              �����    �����    �����              �����    �����    �����              �����    �����    �����              �����    �����    �����              �����    �����    �����              �����                        �����        �����                     ]����       �����       �����                     �����       �����       �����                    �����       �����       �P - �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    ���~��?���  ?����������  ?�~��?���               >0f��3`��  ?����������  ?�~��?���               ?�~��?���  ?����������  ?�~��?���               >0f��3`��  ?����������  ?�~��?���    P ���������                    ������������������������������������          ���������������������������          ���������������������������          ���������������������������                    ���������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z����Wԯ�^�(
P�)@|����>{��������z����Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N��
P�)@|����>{��������r��)�S��)N��
P�)@|����>{��������z��+�Wԯ�^��
P�)@|����>{��������z��+�Wԯ�^��
P�)@|����>{��������s������?�����?�|����>z����Wԯ�^s��)���?���
P�)@|����>z����Wԯ�^s��)���?���
P�)@|����>z����Wԯ�^{��+�������
P�)@|����>z����Wԯ�^{��+�������
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(
P�)@|����>{��������r��)�S��)N�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z��+�W��^�(
P�)@|����>{��������z��+�W��^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(
P�)@|����>{��������r��)�S��)N�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>z��+�W��^s�����?��(
P�)@|����>z��+�W��^s�����?��(
P�)@|����>z��+�W��^{�����ԯ���(
P�)@|����>z��+�W��^{�����ԯ���(
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(
P�)@|����>{��������r��)�S��)N�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(
P�)@|����>{��������r��)�S��)N�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z��+��ԯ�^�(
P�)@|����>{��������z��+��ԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(��)@|����>{��������r��)�S��)N�(��)@|����>{��������z��+�Wԯ�^�(��)@|����>{��������z��+�Wԯ�^�(��)@|����>{��������s������?�����?�|����>z��+��ԯ�^s����S��?��(��)@|����>z��+��ԯ�^s����S��?��(��)@|����>z��+��ԯ�^{����W����(��)@|����>z��+��ԯ�^{����W����(��)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������{��+�W��^�(
P�)@|����>{��������{��+�W��^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(
P�)@|����>{��������r��)�S��)N�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��+�W��^r�����?��(
P�)@|����>{��+�W��^r�����?��(
P�)@|����>{��+�W��^z�����ԯ���(
P�)@|����>{��+�W��^z�����ԯ���(
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ��������������������?���          ������������������~���?�~          ���������x����x����          ���������x����{��������          ���������x����s������?�����?�|����>x����s������?��(
P�)@}k�����_־z��+�Wԯ�^s������?��(
P�)@}k�����_־{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>{��������r��)�S��)N�(
P�)@|����>{��������r��)�S��)N�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������z��+�Wԯ�^�(
P�)@|����>{��������s������?�����?�|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^s������?��(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>z��+�Wԯ�^{���������(
P�)@|����>{��������{������������?�|����>x����x����          ������������������p ���           ���������p ��� p ���           ���������p ��� �����������?����p ��� ������������������          ���������������������������          ���������������������������          ������������������                    ���������                              ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������������������������          ���������?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����