�P  �> P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          UUUUUU   UUUUUU   UUUUUU                       �UUUUU   UUUUUU             �������  �������  �������             ������         �                                �������                       ������         �                                �������                      �������                                         �������                      �������                                        �������                      �������                                        �������                      �������                                    �   �������       �             �������  ���  �  ��  �            ��  �� � ?��� �      @           ���������>  | @                   x   � ��������        >    |  ������}�AD  "��         A    �   wX  � ����O�            ��    ������;�� c��� ��� ��� � @  (� �������� & 2  L d               @ ��������� & 2  L d                 @ ~ ?�0 ~�������                @  � ��  ������  ��  �                 �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P - ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������*���������*���������*���������*���������      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ?���      ?���      ?���      ?���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ��        ��        ��        ��        ��        �        �        �        �        ?�        ?�        ?�        ?�        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �     @�     @�     @�     @�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P  � /�� _ ������  ��    ~ w ?� � ~|  � @>��������  ��     w   � @|w0�`>��������  ��    � �� ��w?���� ����   ���            �w?������������  ��       �    �w?����� ����   ��             �w?�������������  ��             �w?���� ����   ���            �w?���������?���  ���            �w?����� ��0�   ���            �w?���������?���  ���            � ?�� � �����   ����            � ?�� ����������  ��          �  � ?��� � �����   ���        �  � ?��� ����������  ��          �  � ?��� � ��  ��   ��          �  � ?��� ����������  ��  �            � ?��� � ��  ��                     ������������������ ��  ��           ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ �������   �>�    �|>��������|A8 ��   �  8      >��������|�������   �  8      >�������|A�8 ���   �  8      >��������|���������   �  8      >������|A�8?���� ?�� �  8      >��������|��������  � �  8      >��������|A�8 ��  � �  8      >�������|��������  � �  8      ?���������@ 8      �     8      ?����������������?�� ���            �����  �� ��    �             UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ �������   �>�    �|>��������|A8 ��   �  8      >��������|�������   �  8      >�������|A�8 ���   �  8      >��������|���������   �  8      >������|A�8?���� ?�� �  8      >��������|��������  � �  8      >��������|A�8 ��  � �  8      >�������|��������  � �  8      ?���������@ 8      �     8      ?����������������?�� ���            �����  �� ��    �             UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ �������   �>�    �|>��������|A�8 �   �  8      >��������|�������   �  8      >�������|A�8 ��   �  8      >��������|�������   �  8      >������|A8?���� ?�� �  8      >��������|�������   �  8      >��������|A8 ��   �  8      >�������|��������   �  8      ?���������@ 8           8      ?����������������?�� ��            �����  �� ��                 UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ �������   �>�    �|>��������|A�8 �   �  8      >��������|�������   �  8      >�������|A�8 ��   �  8      >��������|�������   �  8      >������|A8?���� ?�� �  8      >��������|�������   �  8      >��������|A8 ��   �  8      >�������|��������   �  8      ?���������@ 8           8      ?����������������?�� ��            �����  �� ��                 UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ ��������   �>�    �|>��������|A�8 ��   �  8      >��������|��������   �  8      >�������|A�8 ���   �  8      >��������|��������   �  8      >������|A8?���� ?�� �  8      >��������|�������  � �  8      >��������|A8 ��  � �  8      >�������|��������  � �  8      ?���������@ 8      �     8      ?����������������?�� ���            �����  �� ��    �             UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ ������   �>�    �|>��������|A8 �   �  8      >��������|������   �  8      >�������|A�8 ��   �  8      >��������|��������   �  8      >������|A�8?���� ?�� �  8      >��������|��������   �  8      >��������|A�8 ��   �  8      >�������|��������   �  8      ?���������@ 8           8      ?����������������?�� ��            �����  �� ��                 UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ ��������   �>�    �|>��������|A�8 ��   �  8      >��������|��������   �  8      >�������|A�8 ���   �  8      >��������|��������   �  8      >������|A8?���� ?�� �  8      >��������|�������  � �  8      >��������|A8 ��  � �  8      >�������|��������  � �  8      ?���������@ 8      �     8      ?����������������?�� ���            �����  �� ��    �             UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                                        ���������                              ���������                      �����  ���������          ?��    ��  �����  ��    ��          ?��    ��  ���  ���������� ?�� �>�    �|  ���  ��?����   �>�����| ������ ������   �>�    �|>��������|A8 �   �  8      >��������|������   �  8      >�������|A�8 ��   �  8      >��������|��������   �  8      >������|A�8?���� ?�� �  8      >��������|��������   �  8      >��������|A�8 ��   �  8      >�������|��������   �  8      ?���������@ 8           8      ?����������������?�� ��            �����  �� ��                 UG��⪨���������   ?��           UG����⪨j���?�UV   �?�           UG����⪨���������                  UG����⪨j��    UV                  UG����⪨���������                  UG����⪨j��    UV                    �����  ���������          UP    
��  �����  ��    ��          UP    
��  �����  ���������                    ���������                              ������������������                    ���������                              ������������������                    ���������                              ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����