�P  `"� M ����������������������������                                                      ���������������������������������������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������                       ���                       ���                           �����������������������������                       ���                       ���                           ��                       ���������������������������������������������������������                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���     � A               �����������������������������                      '����                      '���                     �����������������������������                      '����                      '���                    �����������������������������                      '����                      '���     �O8V8U�Y��       �����������������������������                      '����                      '���     QQDYDUQe$P       �����������������������������                      '����                      '���     �Q|QDUE$P       �����������������������������                      '����                      '���     Q@QDUE$P       �����������������������������                      '����                      '���     $QQD�D�QE$P       �����������������������������                      '����                      '���     ÎO8�8��D��       �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���        @            �����������������������������                      '����                      '���         @            �����������������������������                      '����                      '���         @            �����������������������������                      '����                      '���     J���5N�<�,        �����������������������������                      '����                      '���     K*,�(�A YD(�        �����������������������������                      '����                      '���     �*�(�O�D/�        �����������������������������                      '����                      '���     �*�(�QQD("        �����������������������������                      '����                      '���     *(�(�QQD(�        �����������������������������                      '����                      '���     )ȁ�%O�<
'"�       �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���         �                �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ����������������  ����������             ���     '����                      '���      y@@  �   ���        �����������������������������             ���     '����             ���     '���      � @ �   ���        ����������������  ����������                    '����                    '���      � @ �   ���        ���������������� ����������                    '����                    '���      �NH��ǫ ���        ���������������� ����������                    '����                    '���      �QP �(�����        ����������������?�����������                    '����                    '���      �P` �言��        ����������������?�����������                    '����                    '���      �PP �����        ����������������?�����������                    '����                    '���      �QH �(����        ���������������� ����������                    '����                    '���      yND	��Ǩ����        ���������������� ����������                    '����                    '���             � ���        ����������������  ����������                    '����                    '���              ���        ����������������  ����������             ���     '����             ���     '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ��                       ���������������������������������������������������������                           �����������������������������                       ���                       ���                           �����������������������������                       ���                       ���                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                                                       ��������������������������������������������������������                                          (�(                            ( �� Q8Q��@�Or'�@���D�E� ������������������������������ �(                            (�(                          