�P  �]�8                                                                                                                                                                                                                                                              �            �           �             �                    ��           �                         @                                x           �             �                                                                             �  ��           �           �             �                �                                                           �  ?��           �           �             �                                                                             ��� ��          �           �             �               �                                                          �� ��           �           �             �                                                                            ������          ��          �             �                                                                           ��� ���          �           �             �                                                                            ���/���          �           �             �                                                                          ������          ��          �             �                                                                            �������     �� ��� ~� ?�8 �        � p �     � � �               �   @ � � �D            �        �    �������     �� ��� ~  �8 �        � p �     �� �                                                                �������     ������ ������ �        ��� �    ���� ��                  @    �              @           � @ ?�������     ������ �?���| �        ��� �    ��� ��                                                               ?�������    ������������� �        ��� �    ?�������� @                        	                             �    ?�������     �������������� �        ?��� �    �������                                                               �������    �����������������        ���� �    ?��������                                            
                  �������    �������������� �        ��� �    ��������                                                               �������    ��������������� ��x   ���� �   ���������                 @                 �                        �������    �����������������  �    ���� �    ���������                                                               �������    ����� ��������������   ���� �  ���������                                                             �������    �����������������?��   ���� �  ���������                                                               �������    ����� ��������������   ������ ����������                                                            �������    ����� ��������������   ���� � ����������                                                               �������    ?����� ��������������   ���� � ����������                                                  @          �������    ����� ��������������   ������ ?����������                                                               ������@ � ?����� ��������������   ������ ����������                                                          ������� � ?����� ��������������   ������ ����������                                                               ������  ��@?����� ���������������  �����������������                                 � �                        ������  ���?����� ��������������   ������ �����������                                                               ?������ ���?����� ��?�������������  �����������������                   �                                      ������ ���?����� ��?�������������  �����������������                                                               ����� ���?����� ����������������  ����������������� @ $                 �                                    ?���~� ���?����� ���������������  �����������������                                                               �� ?� ?���?����� ����������������  ?�����������������                                     @                        ?�� � ���?����� ����������������  �����������������                                                               ?�� � ?�������� ����������������  ?�����������������     @  @                                                 ?�� ?� ?�������� ����������������  ?�����������������                                                               ?�?� � �������� ����������������  ?����������������        �          @     @         @                 ?�� ?� �������� ����������������  ?�����������������                                                               ?��� ?���������� ������� ����?��  ����������� _�                       @                     �                ?��� ?� ��������� ���� �  ��������  ��}��������� ?�                                                                 ?��� ?���������� �����  ?  ��������  � =��������� �                    �                      @              ?��� ?���������� ����    �������  � ��������� �                                                                 ?��� ?����������������  ?  ��?������  �� ����� ���� �                                       �    @              ?��� ?���������������  ?  �������  � ��?������� �                                                                 ?��� ?�����������������    ��������  �� ���������� �                                                               ?��� ?�����������������    ���������  �� ������ ���� �                                                                 ?��� �����������������    ���������  �� ����������� �                             �                      �         ?��� ?����������������    ���������  �� ������ ���� �                                                                 ?��� ����������������  ?� ��������� �� ����������� �        @          �         �                                ?��� ?���������������    ���������  �� ����������� �                                                                 ?��� ?���������������  ?� ���������  �� ����������� �                              �                      @        ?��� ���������������    ��������� �� ����������� �                                                                 ?��� ���������������  ?  ��������� �  ����?������� �                        � @                                   ?��� ��������������  ?� ��������� �� ����������� �                                                                 ?��� ���������������  ?� �������� �   ����?������� �               ( �                                    !         ?��� ��������������  ?� ��������� �  ����?������� �                                                                 ��� �������������?��  � ��������� �  ����������� �                                                                 ?��� ��������������   ?� ��������� �  ����?������  �                                                                 ?��� ��������������   � ��������� �  �����������  �                                                @            ��� �������������?�   � ��������� � �����?������  �                                                                 ?��� �������������?�   �� ��������� � �����������  �                                                                ��� ������������?�   � ��������� � �����������  �                                                                 ��� ������������?�   � �������� � ������������ �                                     @                       ��� �������������   �� ��������� � �����������  �                                                                 ��� �������������  �� �������� � ������������ �                                            �     @      ��� �������������   �� �������� � ������������ �                                                                 ��� �������������   �� ������ � ������������� �                 �          @                            ��� �������������  �� ������� � ������������� �                                                                 �������������������  �� �����<� � ������������� �         @        @         @      @                       ������� ����������  �� ?�����>� � ?������������ �                                                                 ���?���� ����������  �� ����� � � ?�?���������� ?�                                                          ������� ��������?��  �� ?���� � � ����������� �                                                                 �������� ��������?��  �� ���� �  ���?���������� ?�       �                                               `        ������� ������� ?��  �� ���� � ����?���������� ?�                                                                 �������� ������ ?��  �� ���� � ����?��������� �                                               H            �������� ���?��� ?��  �� ���� �  �������������� ?�                                                                 �������� �������?��  �� ���� �  �������������� ?�                                                             �������� ������ ?��  �� ���� �  ������������� �                                                                 ��������������� ?��  �� ���� �  ��������?���� �                                                   @           �����������������?��  �� ���� �  �������?�� �� �                                                                 �����������������?��  �� ���� �  ?��������� ?� �                                               �            �����������������?��  �� ���� �  ������ �� � �                                                                 ������������� ����?��  �� ���� �  ?��������� � �                    @                                       ������������� ����?��  �� ���� �  ?������ �� � �                                                                 ������������� ����?��  �� ���� �  ?������ �� � �             @                                              ������������� ���?��  �� ���� �  ������ �� � �                                                                  ������������ ���?��  �� ���� �  ������  �� � �                                                             ������������� ?�����  �� � ��� �  ������  �� � �                                                                  ������������ ����  �� � ���  �  ������  �� � ?�                                 �               �          ���������� �����  �� � ��  �  ���� ��  � � �                                                                  ?�����?���� �����  �� � ��  �  ���� ��  ~�  x �                     @          @          @  �               � ?������� ����  �� � ?��  �  ���� �  �  � ?�                                                                  � ��|���� �?���  �� � ?�  ~  �� � �  ~�  x ?�              �@             �   �           @   8       � �������   ?���  �� � �  ~   �� � ?�  >�    �                                                                     �� ����   � ��   �  � �  >   � � �  |�    �        �$ �               �@       @                        �  ���     ��   �  � �  <   � � �  >~    �                                                                                      �          �            �                                                                                                �          �             �                                                                                                �          �             �                                                                                                �          �             |                                                                                                p          �                                                           @                                                  �          ?�                                                                                                                         ?�                                                                                                                          ?�                                                                                                                          �                                                                                                                          �                                                                                                                                                                                                                                                                                                                                                                                                                                                             Y                                                                        �                                                                                                                                                      �                                                                                  0  �                 |             �                      �      ���                          @             �                      �      �       `  �                 >             |                      |    � |�                                                                                 0v??�� �       �   ;��   p       �w��8���         �w� �������      @� �        �  %    H        J$	R�  �       J �
       w?�� `       �   ��  0 0       �1����|         �1� ������                                                                               ��w����� x       ��@ ?��  < <       �����������      �����������    �              @      @             �   � @          Q    @    8w���� �       ��  ?��  8 x       ���<�����      ����������                                                                               ��w������� �     �X` ?�� x`| >     ��������������    ��������� �   �  ` �         $�    D@        �   �     $ @       �  �       ��w?����`� �     ��p ?�� 80x >     ���<�������    ��������� �                                                                             ��s����     �p�?��_�|�� A     �����|�o��    ����߾��Ϟ��    @   A              �          �D �  �@�       �@  @@  �   ��w��ߏ���     �<�~��?8px A     ��?��<�>������    ��?���?���� �            �                   >                                          � ��w��ß���     �?���8����� ��     s���|�|1���π     s��ώ�s� �                    �   @                         �             @    ��s��Ï��     �>���8�<�x ��     s烃�<�<`���     s烇ߎ�qϜ �           �                                                            � ��y������     ן����9����� @     s���x�x ���      s��ߎ�p��x�               �       ! �           !D !@  0��        �   0   �����Î��     �?����8�ߜ�p @     s��8�8 ���� �     s���qϞ��           �                   ��                                        � ����o�����     ������8����� @     q������ ����      q�����p�?��  
  @              @      �            @       �             �    ��������     ������9����p @     s����8�p ���� �     s�����p���           �                   ��                                        � ����ǜ���     ������y����p @     �����������      �������?��                 @                    �  �     �        @         ����Ü��     ������9����� @     q����p�p ���� �     q�����p���           �                   ��                                        � ������s���     ������=����` @     {߇����������      {߇���x���               @  @	          �   �   �     �     �    ��   �����Ü;��     �����9����� @     q߃��p�p����� �     q߃���p~>�           �                   ��                                        � ����������     �8?�����=��� @     �ǃ�����������     �ǃ��À��`�   �   �           $@                  &   &     �        �   0   �8������     �8�������� @    �χ��s���y�����x�    �χ��?���~> �           �                   ��                                        � p9�����_��     ��=�����������    �Ç�������������    �Ç������~?��     @  �                   @                 @     �                   �8�����?��     �������������    �Ç�����?�������    �Ç���Ǉ�|?��           �                                                            � �9��������     �����������A     ������������c��    �����ǃ�<?�� �   �               @                            �                 `8��?����     �����������A     ����������������    ������Ǉ�x?��            �                   >                                          � p1����� �     �����?�x >     ���������?�7��    �����ǁ�p?� �    �            �   H  �          B�    @             @     `�~��� �     �������x >     ����������~�7��    ������Ã�8� �                                                                                @             �       �                    x             �     X      �                      �                                                 `             �                     �  �   �             �     <                                                                                                                                                                                                                                                         8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                                                                                                                                                                                                                                                                                                  �      �  �` Ϙ<y�` > �                                                                                                    �          `���3f�` 3 �3                                                                                                     �           `��f�0` 3 �0                                                                                                     ��m�s���ݟ|�f�0|l3<�0<}�|                                                                                                 ���m�f`6fٳv��f�`fl>f�f͛v                                                                                                 ����g��6fٳf��f�`fl3f�~͛f                                                                 ��0�f 6fٳf��f��fl3f�`͛f                                                                                                 ���33f`6c��f���0f��f83f�3fͻf                                                                                                 ��3c�����fa��?<x�|0><�<|�f                                                                                                            �     0                                                                                                                  >  �     �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �                                                                                            �                                                             ������     �                                                       ͍�6f                                                            ͍��                                                            ͍��q������                                                    ������ٶ�0lٳ��                                                   ͍�6l�a��3��3�                                  ͍�6f 1��6l�3�                                                   ͍�6� ���6lٳـ                                                   �������p�����g��                                                           �                                                                 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  