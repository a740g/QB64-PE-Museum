�P  `"� M ����������������������������                                                      ���������������������������������������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������                       ���                       ���                           �����������������������������                       ���                       ���                           ��                       ���������������������������������������������������������                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���            �           �����������������������������                      '����                      '���             �            �����������������������������                      '����                      '���        @    �            �����������������������������                      '����                      '���        �"��`          �����������������������������                      '����                      '���        ��R���          �����������������������������                      '����                      '���        ��R��@          �����������������������������                      '����                      '���        ��R��           �����������������������������                      '����                      '���        ��R���          �����������������������������                      '����                      '���        �󒧂`          �����������������������������                      '����                      '���                          �����������������������������                      '����                      '���           �              �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������    `` �  �  8    '����    `` �  �  8    '���      `` �  �  8       �����������������������������   ��� �����    '����   ��� �����    '���     ��� �����       �����������������������������   �?�� ����    '����   �?�� ����    '���     �?�� ����       ��������?����������w���������   �?�<?� �ǻ���    '����   �<8<;� �ǁ��p    '���     �?�<?� �ǻ���       ��������?�������~7���������   �?�<� �������    '����   �<<8q� ��Ǉ0    '���     �?�<� �������       ����������������|����������   �|~|���ρ�ϟp    '����   �|~p� ����     '���     �|~|���ρ�ϟp       ����������������������������   �<~�������>>    '����   �~��p����8    '���     �<~�������>>       ��������������>�������������   �|s������|    '����   �8c����x    '���     �|s������|       ������@� ?  !�@�����������      @ � �     '����                      '���     �9���������x       ������� >� ��������������    �  @       '����                      '���     �8������x>       �������x  �������������    �	   � $      '����                      '���     �y�����=�p�       �������p� a������������      (          '����                      '���     �<�����>�q�       �������0<`� `�����������    `@    � d    '����                      '���     �x�ß�����s�       ������ �8< ?� G�����������   � 78 �@�    '����                      '���     �}�����߸8��       ������`><b?� �ǌG���������   �@C�@��s�    '����                      '���     ���Ý����88s�       ��������?>?�?0�������������   q���@�π8?    '����                      '���     q�����π8?8       �������~������������������    ��  ` 00 0    '����                      '���      ��  ` 00 0       ����������������������������        �       0    '����                      '���          �       0       �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ����������������  ����������             ���     '����                      '���      y@@  �   ���        �����������������������������             ���     '����             ���     '���      � @ �   ���        ����������������  ����������                    '����                    '���      � @ �   ���        ���������������� ����������                    '����                    '���      �NH��ǫ ���        ���������������� ����������                    '����                    '���      �QP �(�����        ����������������?�����������                    '����                    '���      �P` �言��        ����������������?�����������                    '����                    '���      �PP �����        ����������������?�����������                    '����                    '���      �QH �(����        ���������������� ����������                    '����                    '���      yND	��Ǩ����        ���������������� ����������                    '����                    '���             � ���        ����������������  ����������                    '����                    '���              ���        ����������������  ����������             ���     '����             ���     '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           �����������������������������                      '����                      '���                           ��                       ���������������������������������������������������������                           �����������������������������                       ���                       ���                           �����������������������������                       ���                       ���                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                           �����������������������������������������������������������������������������������                                                       ��������������������������������������������������������                                          (�(                            ( �� Q8Q��@�Or'�@���D�E� ������������������������������ �(                            (�(                          