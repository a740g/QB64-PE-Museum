�P  �> P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������                  �������  �������  �������  �������  ffffff`  �������  9�������  9�������  ffffff`  �������  �������  �������  &ffffffd  �������  �������  �������  &ffffffd  �������  �������  �������  &ffffffd  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  &d  �������  �������  �������  ffffffd ���������                  ���������	���������	���������	���������ffffffff`���������������������������ffffffff ���������������������������$ffffffff$���������������������������dffffffff&���������������������������dffffffff&���������������������������dffffffff&���������������������������dffffffff&���������������������������dffffffff&     �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P - ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ���      ��        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P ���������        X        Xe������������������������������������ffffffffff���������������������������ffffffffff����������      	��      	�fo�������f�      	��      	��      	�fo�������f�      	��      	��      	�fo�������f�      	��      	��      	�fo�������f�9�q�	��      	��      	�fo�s�0��f�R�(�	��      	��      	�fo��w�]�f�=ȁ�	��      	��      	�fo��7~A�f�E�(�	��      	��      	�fo���}�_�f�ER�(�	��      	��      	�fo��u�]�f�=�q�	��      	��      	�fo�s���f�    	��      	��      	�fo�������f�    	��      	��      	�fo�������f�      	��      	��      	�fo�������f�      	��      	��      	�fo�������f�      	�������������������f`      f���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff � � � � � �g��������~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f�~����~�� � � � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � ��~����~�� � �f�`h�`f � � � � � �g������� � � � � � �g������� � � � � � �g������� � � � � � �g����������������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff���������������������������ffffffffff?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����